VERSION 5.4 ;
NAMESCASESENSITIVE ON ;

UNITS
    DATABASE MICRONS 1000  ;
END UNITS

LAYER PC
    TYPE MASTERSLICE ;
END PC

LAYER CA
    TYPE CUT ;
END CA

LAYER metal1
    TYPE ROUTING ;
    WIDTH 0.160 ;
	AREA 0.089 ;
    SPACING 0.160 ;
    SPACING .26 RANGE 1.77 4.00 ;
    SPACING .36 RANGE 4.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.400 ;
    DIRECTION HORIZONTAL ;
	MINIMUMCUT 2 WIDTH 1.04 ;
    RESISTANCE RPERSQ 0.07090000 ;
	CAPACITANCE CPERSQDIST 9.7045e-05 ;
	EDGECAPACITANCE 8.3040e-05 ;
END metal1

LAYER V1
    TYPE CUT ;
	SPACING 0.28 ;
END V1

LAYER metal2
    TYPE ROUTING ;
    WIDTH 0.200 ;
	AREA 0.120 ;
    SPACING 0.200 ;
    SPACING .28 RANGE 2.01 4.00 ;
    SPACING .36 RANGE 4.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.400 ;
    DIRECTION VERTICAL ;
	MINIMUMCUT 2 WIDTH 1.04 ;
    RESISTANCE RPERSQ 0.06390000 ;
	CAPACITANCE CPERSQDIST 9.9389e-05 ;
	EDGECAPACITANCE 7.1337e-05 ;
END metal2

LAYER V2
    TYPE CUT ;
	SPACING 0.28 ;
END V2

LAYER metal3
    TYPE ROUTING ;
    WIDTH 0.200 ;
	AREA 0.120 ;
    SPACING 0.200 ;
    SPACING .28 RANGE 2.01 4.00 ;
    SPACING .36 RANGE 4.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.400 ;
    DIRECTION HORIZONTAL ;
	MINIMUMCUT 2 WIDTH 1.04 ;
    RESISTANCE RPERSQ 0.06390000 ;
	CAPACITANCE CPERSQDIST 9.1182e-05 ;
	EDGECAPACITANCE 7.1611e-05 ;
END metal3

LAYER V3
    TYPE CUT ;
	SPACING 0.28 ;
END V3

LAYER metal4
    TYPE ROUTING ;
    WIDTH 0.200 ;
	AREA 0.120 ;
    SPACING 0.200 ;
    SPACING .28 RANGE 2.01 4.00 ;
    SPACING .36 RANGE 4.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.400 ;
    DIRECTION VERTICAL ;
	MINIMUMCUT 2 WIDTH 1.04 ;
    RESISTANCE RPERSQ 0.06390000 ;
	CAPACITANCE CPERSQDIST 8.4534e-05 ;
	EDGECAPACITANCE 7.1142e-05 ;
END metal4

LAYER VL
    TYPE CUT ;
	SPACING 0.56 ;
END VL

LAYER metal5
    TYPE ROUTING ;
    WIDTH 0.400 ;
	AREA 0.480 ;
    SPACING 0.400 ;
    SPACING .60 RANGE 2.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.800 ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.03730000 ;
	CAPACITANCE CPERSQDIST 6.6102e-05 ;
	EDGECAPACITANCE 7.1227e-05 ;
END metal5

LAYER VQ
    TYPE CUT ;
	SPACING 0.56 ;
END VQ

LAYER metal6
    TYPE ROUTING ;
    WIDTH 0.400 ;
	AREA 0.480 ;
    SPACING 0.400 ;
    SPACING .60 RANGE 2.01 8.00 ;
    SPACING 1.12 RANGE 8.01 25.00 ;
    SPACING 1.92 RANGE 25.01 100000.0 ;
    PITCH 0.800 ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.03730000 ;
	CAPACITANCE CPERSQDIST 3.5152e-05 ;
	EDGECAPACITANCE 6.8060e-05 ;
END metal6

VIA via1 DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal1 ;
        RECT -0.120 -0.160 0.120 0.160 ;
    LAYER V1 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via1

VIA via1r DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal1 ;
        RECT -0.160 -0.120 0.160 0.120 ;
    LAYER V1 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via1r

VIA via1_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal1 ;
        RECT -0.120 -0.360 0.120 0.360 ;
    LAYER V1 ;
        RECT -0.100 0.100 0.100 0.300 ;
        RECT -0.100 -0.300 0.100 -0.100 ;
    LAYER metal2 ;
        RECT -0.100 -0.300 0.100 0.300 ;
END via1_fat

VIA via1r_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal1 ;
        RECT -0.360 -0.120 0.360 0.120 ;
    LAYER V1 ;
        RECT -0.300 -0.100 -0.100 0.100 ;
        RECT 0.100 -0.100 0.300 0.100 ;
    LAYER metal2 ;
        RECT -0.300 -0.100 0.300 0.100 ;
END via1r_fat

VIA via2 DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER V2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via2

VIA via2ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 6.000 ;
    LAYER metal2 ;
        RECT -0.100 -0.300 0.100 0.300 ;
    LAYER V2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via2ts

VIA via2_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal2 ;
        RECT -0.100 -0.300 0.100 0.300 ;
    LAYER V2 ;
        RECT -0.100 0.100 0.100 0.300 ;
        RECT -0.100 -0.300 0.100 -0.100 ;
    LAYER metal3 ;
        RECT -0.100 -0.300 0.100 0.300 ;
END via2_fat

VIA via2r_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal2 ;
        RECT -0.300 -0.100 0.300 0.100 ;
    LAYER V2 ;
        RECT -0.300 -0.100 -0.100 0.100 ;
        RECT 0.100 -0.100 0.300 0.100 ;
    LAYER metal3 ;
        RECT -0.300 -0.100 0.300 0.100 ;
END via2r_fat

VIA via3 DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER V3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal4 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via3

VIA via3ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 6.000 ;
    LAYER metal3 ;
        RECT -0.300 -0.100 0.300 0.100 ;
    LAYER V3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
    LAYER metal4 ;
        RECT -0.100 -0.100 0.100 0.100 ;
END via3ts

VIA via3_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal3 ;
        RECT -0.100 -0.300 0.100 0.300 ;
    LAYER V3 ;
        RECT -0.100 0.100 0.100 0.300 ;
        RECT -0.100 -0.300 0.100 -0.100 ;
    LAYER metal4 ;
        RECT -0.100 -0.300 0.100 0.300 ;
END via3_fat

VIA via3r_fat DEFAULT
    RESISTANCE 6.000 ;
    LAYER metal3 ;
        RECT -0.300 -0.100 0.300 0.100 ;
    LAYER V3 ;
        RECT -0.300 -0.100 -0.100 0.100 ;
        RECT 0.100 -0.100 0.300 0.100 ;
    LAYER metal4 ;
        RECT -0.300 -0.100 0.300 0.100 ;
END via3r_fat

VIA via4 DEFAULT
    RESISTANCE 3.000 ;
    LAYER metal4 ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER VL ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER metal5 ;
        RECT -0.200 -0.200 0.200 0.200 ;
END via4

VIA via4ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 3.000 ;
    LAYER metal4 ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER VL ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER metal5 ;
        RECT -0.200 -0.200 0.200 0.200 ;
END via4ts

VIA via5 DEFAULT
    RESISTANCE 3.000 ;
    LAYER metal5 ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER VQ ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER metal6 ;
        RECT -0.200 -0.200 0.200 0.200 ;
END via5

VIA via5ts DEFAULT TOPOFSTACKONLY
    RESISTANCE 3.000 ;
    LAYER metal5 ;
        RECT -0.600 -0.200 0.600 0.200 ;
    LAYER VQ ;
        RECT -0.200 -0.200 0.200 0.200 ;
    LAYER metal6 ;
        RECT -0.200 -0.200 0.200 0.200 ;
END via5ts

VIARULE via1Array GENERATE
    LAYER metal1 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.060 ;
        METALOVERHANG 0.000 ;

    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER V1 ;
        RECT -0.100 -0.100 0.100 0.100 ;
        SPACING 0.600 BY 0.600 ;
END via1Array

VIARULE via2Array GENERATE
    LAYER metal2 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER V2 ;
        RECT -0.100 -0.100 0.100 0.100 ;
        SPACING 0.600 BY 0.600 ;
END via2Array

VIARULE via3Array GENERATE
    LAYER metal3 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER V3 ;
        RECT -0.100 -0.100 0.100 0.100 ;
        SPACING 0.600 BY 0.600 ;
END via3Array

VIARULE via4Array GENERATE
    LAYER metal4 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER VL ;
        RECT -0.200 -0.200 0.200 0.200 ;
        SPACING 0.800 BY 0.800 ;
END via4Array

VIARULE via5Array GENERATE
    LAYER metal5 ;
        DIRECTION HORIZONTAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER metal6 ;
        DIRECTION VERTICAL ;
        OVERHANG 0.000 ;
        METALOVERHANG 0.000 ;

    LAYER VQ ;
        RECT -0.200 -0.200 0.200 0.200 ;
        SPACING 0.800 BY 0.800 ;
END via5Array

VIARULE TURNmetal1 GENERATE
    LAYER metal1 ;
        DIRECTION vertical ;

    LAYER metal1 ;
        DIRECTION horizontal ;
END TURNmetal1

VIARULE TURNmetal2 GENERATE
    LAYER metal2 ;
        DIRECTION vertical ;

    LAYER metal2 ;
        DIRECTION horizontal ;
END TURNmetal2

VIARULE TURNmetal3 GENERATE
    LAYER metal3 ;
        DIRECTION vertical ;

    LAYER metal3 ;
        DIRECTION horizontal ;
END TURNmetal3

VIARULE TURNmetal4 GENERATE
    LAYER metal4 ;
        DIRECTION vertical ;

    LAYER metal4 ;
        DIRECTION horizontal ;
END TURNmetal4

VIARULE TURNM5 GENERATE
    LAYER metal5 ;
        DIRECTION vertical ;

    LAYER metal5 ;
        DIRECTION horizontal ;
END TURNM5

VIARULE TURNM6 GENERATE
    LAYER metal6 ;
        DIRECTION vertical ;

    LAYER metal6 ;
        DIRECTION horizontal ;
END TURNM6

SPACING
    SAMENET metal1 metal1 0.160  ;
    SAMENET metal2 metal2 0.200 STACK ;
    SAMENET metal3 metal3 0.200 STACK ;
    SAMENET metal4 metal4 0.200 STACK ;
    SAMENET metal5 metal5 0.400 STACK ;
    SAMENET metal6 metal6 0.400  ;
    SAMENET V1 V1 0.200  ;
    SAMENET V2 V2 0.200  ;
    SAMENET V3 V3 0.200  ;
    SAMENET VL VL 0.400  ;
    SAMENET VQ VQ 0.400  ;
    SAMENET V1 V2 0.0 STACK ;
    SAMENET V2 V3 0.0 STACK ;
    SAMENET V3 VL 0.0 STACK ;
    SAMENET VL VQ 0.0 STACK ;
END SPACING

SITE cellsite
    SYMMETRY y  ;
    CLASS core  ;
    SIZE 0.400 BY 3.600 ;
END cellsite

MACRO MAS1
    CLASS CORE ;
    FOREIGN MAS1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.360 0.920 1.520 3.160 ;
        RECT  0.920 0.920 1.360 1.080 ;
        RECT  1.280 1.910 1.360 3.160 ;
        RECT  1.040 1.910 1.280 2.750 ;
        RECT  0.640 0.800 0.920 1.080 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.430 0.680 1.710 ;
        RECT  0.320 1.240 0.360 1.710 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.240 1.160 1.700 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.470 -0.280 1.600 0.280 ;
        RECT  1.160 -0.280 1.470 0.760 ;
        RECT  0.450 -0.280 1.160 0.280 ;
        RECT  0.150 -0.280 0.450 1.080 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.520 3.320 1.600 3.880 ;
        RECT  0.240 2.530 0.520 3.880 ;
        RECT  0.000 3.320 0.240 3.880 ;
        END
    END VDD
END MAS1

MACRO MAS10
    CLASS CORE ;
    FOREIGN MAS10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.350 0.840 1.520 2.940 ;
        RECT  1.280 0.840 1.350 1.960 ;
        RECT  1.230 2.230 1.350 2.940 ;
        RECT  1.200 0.840 1.280 1.220 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.680 1.240 0.720 1.560 ;
        RECT  0.480 1.240 0.680 1.750 ;
        RECT  0.400 1.470 0.480 1.750 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.000 -0.280 1.600 0.280 ;
        RECT  0.720 -0.280 1.000 1.080 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.030 3.320 1.600 3.880 ;
        RECT  0.750 2.230 1.030 3.880 ;
        RECT  0.000 3.320 0.750 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  0.950 1.520 1.120 2.070 ;
        RECT  0.530 1.910 0.950 2.070 ;
        RECT  0.240 1.910 0.530 2.350 ;
        RECT  0.240 1.030 0.320 1.310 ;
        RECT  0.230 1.030 0.240 2.350 ;
        RECT  0.080 1.030 0.230 2.070 ;
    END
END MAS10

MACRO MAS11
    CLASS CORE ;
    FOREIGN MAS11 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.000 1.240 1.120 2.360 ;
        RECT  0.960 0.440 1.000 2.360 ;
        RECT  0.840 0.440 0.960 3.160 ;
        RECT  0.680 0.440 0.840 1.310 ;
        RECT  0.680 1.910 0.840 3.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 1.470 0.680 1.750 ;
        RECT  0.360 1.240 0.400 1.750 ;
        RECT  0.080 1.240 0.360 2.360 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 -0.280 1.200 0.280 ;
        RECT  0.160 -0.280 0.440 0.990 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 3.320 1.200 3.880 ;
        RECT  0.160 2.750 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
END MAS11

MACRO MAS12
    CLASS CORE ;
    FOREIGN MAS12 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.610 6.050 1.520 ;
        RECT  4.810 0.610 5.890 0.770 ;
        RECT  4.650 0.610 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.150 1.640 8.320 2.390 ;
        RECT  7.980 1.030 8.150 2.390 ;
        RECT  7.870 1.030 7.980 1.310 ;
        RECT  7.870 2.110 7.980 2.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.880 0.470 9.120 3.140 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.630 -0.280 9.200 0.280 ;
        RECT  8.350 -0.280 8.630 1.220 ;
        RECT  6.490 -0.280 8.350 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.630 3.320 9.200 3.880 ;
        RECT  8.350 2.990 8.630 3.880 ;
        RECT  7.380 3.320 8.350 3.880 ;
        RECT  7.100 3.260 7.380 3.880 ;
        RECT  6.250 3.320 7.100 3.880 ;
        RECT  5.800 3.200 6.250 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  8.560 1.590 8.720 2.710 ;
        RECT  7.230 2.550 8.560 2.710 ;
        RECT  7.670 0.450 7.810 0.670 ;
        RECT  7.690 1.670 7.760 1.950 ;
        RECT  7.670 1.670 7.690 2.350 ;
        RECT  7.510 0.450 7.670 2.350 ;
        RECT  7.410 2.070 7.510 2.350 ;
        RECT  7.230 1.030 7.350 1.250 ;
        RECT  7.070 1.030 7.230 2.710 ;
        RECT  6.290 1.900 7.070 2.060 ;
        RECT  6.490 2.430 7.070 2.710 ;
        RECT  6.660 2.870 6.940 3.140 ;
        RECT  5.730 2.870 6.660 3.030 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 1.020 5.730 3.030 ;
        RECT  5.450 1.020 5.570 1.310 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.890 1.170 5.170 1.830 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.890 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.590 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END MAS12

MACRO MAS13
    CLASS CORE ;
    FOREIGN MAS13 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 0.780 2.150 2.760 ;
        RECT  1.760 0.780 1.990 1.060 ;
        RECT  1.680 2.440 1.990 2.760 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.520 2.940 2.290 3.100 ;
        RECT  1.280 2.770 1.520 3.160 ;
        RECT  0.570 2.770 1.280 2.930 ;
        RECT  0.260 2.650 0.570 2.930 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.860 1.100 2.140 ;
        RECT  0.480 1.860 0.760 2.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.860 1.190 3.120 2.360 ;
        RECT  2.630 1.190 2.860 1.630 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.010 -0.280 3.200 0.280 ;
        RECT  2.730 -0.280 3.010 1.030 ;
        RECT  1.020 -0.280 2.730 0.340 ;
        RECT  0.720 -0.280 1.020 1.030 ;
        RECT  0.000 -0.280 0.720 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.000 3.320 3.200 3.880 ;
        RECT  2.720 2.550 3.000 3.880 ;
        RECT  0.970 3.320 2.720 3.880 ;
        RECT  0.660 3.200 0.970 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.310 0.930 2.470 2.780 ;
        RECT  1.670 1.220 1.830 2.200 ;
        RECT  1.560 1.220 1.670 1.380 ;
        RECT  1.490 2.040 1.670 2.200 ;
        RECT  1.280 0.930 1.560 1.380 ;
        RECT  1.270 1.540 1.510 1.880 ;
        RECT  1.300 2.040 1.490 2.490 ;
        RECT  0.370 1.540 1.270 1.700 ;
        RECT  0.320 0.930 0.370 1.700 ;
        RECT  0.160 0.930 0.320 2.490 ;
        RECT  0.090 0.930 0.160 1.210 ;
        RECT  0.090 2.210 0.160 2.490 ;
    END
END MAS13

MACRO MAS14
    CLASS CORE ;
    FOREIGN MAS14 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 0.440 2.320 2.720 ;
        RECT  2.080 0.440 2.160 1.560 ;
        RECT  1.760 2.440 2.160 2.720 ;
        RECT  1.390 0.900 2.080 1.060 ;
        RECT  1.110 0.780 1.390 1.060 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.220 1.120 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.220 1.560 1.570 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 1.240 0.720 1.560 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.790 -0.280 2.400 0.280 ;
        RECT  0.590 -0.280 1.790 0.340 ;
        RECT  0.000 -0.280 0.590 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 3.320 2.400 3.880 ;
        RECT  0.600 2.800 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.880 1.580 1.920 1.860 ;
        RECT  1.720 1.580 1.880 2.280 ;
        RECT  0.370 2.120 1.720 2.280 ;
        RECT  0.240 0.800 0.370 1.080 ;
        RECT  0.240 1.920 0.370 2.280 ;
        RECT  0.080 0.800 0.240 2.280 ;
    END
END MAS14

MACRO MAS15
    CLASS CORE ;
    FOREIGN MAS15 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 0.900 2.720 2.800 ;
        RECT  2.410 0.900 2.480 1.140 ;
        RECT  1.910 2.520 2.480 2.800 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.520 1.200 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 2.030 2.070 2.360 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.220 2.700 1.540 3.160 ;
        RECT  0.760 2.700 1.220 2.880 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.370 0.410 1.650 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.140 -0.280 2.800 0.280 ;
        RECT  1.460 -0.280 2.140 0.340 ;
        RECT  0.410 -0.280 1.460 0.280 ;
        RECT  0.130 -0.280 0.410 0.460 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.420 3.320 2.800 3.880 ;
        RECT  2.140 3.200 2.420 3.880 ;
        RECT  0.410 3.320 2.140 3.880 ;
        RECT  0.130 2.800 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.040 1.580 2.260 1.870 ;
        RECT  1.970 0.660 2.190 1.250 ;
        RECT  1.520 1.580 2.040 1.740 ;
        RECT  1.220 0.660 1.970 0.820 ;
        RECT  1.360 1.170 1.520 2.400 ;
        RECT  1.170 1.170 1.360 1.330 ;
        RECT  0.860 2.240 1.360 2.400 ;
        RECT  0.930 0.540 1.220 0.820 ;
        RECT  0.890 1.010 1.170 1.330 ;
        RECT  0.580 2.210 0.860 2.490 ;
    END
END MAS15

MACRO MAS16
    CLASS CORE ;
    FOREIGN MAS16 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.040 0.840 3.120 1.960 ;
        RECT  2.880 0.840 3.040 2.680 ;
        RECT  2.870 1.000 2.880 1.280 ;
        RECT  1.640 2.520 2.880 2.680 ;
        RECT  2.110 1.120 2.870 1.280 ;
        RECT  1.950 1.000 2.110 1.280 ;
        RECT  1.380 2.380 1.640 2.680 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.620 1.010 1.780 ;
        RECT  0.480 1.620 0.720 1.980 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.190 1.760 1.350 2.100 ;
        RECT  1.120 1.940 1.190 2.100 ;
        RECT  0.880 1.940 1.120 2.360 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.560 2.720 2.040 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 1.440 2.320 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.600 1.640 1.920 2.040 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 -0.280 3.200 0.280 ;
        RECT  0.950 -0.280 1.280 1.190 ;
        RECT  0.370 -0.280 0.950 0.280 ;
        RECT  0.090 -0.280 0.370 0.600 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.850 3.320 3.200 3.880 ;
        RECT  2.570 2.840 2.850 3.880 ;
        RECT  0.430 3.320 2.570 3.880 ;
        RECT  0.270 2.520 0.430 3.880 ;
        RECT  0.000 3.320 0.270 3.880 ;
        END
    END VDD
END MAS16

MACRO MAS17
    CLASS CORE ;
    FOREIGN MAS17 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.850 1.920 3.160 ;
        RECT  1.200 0.850 1.760 1.130 ;
        RECT  1.600 1.940 1.760 3.160 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.610 1.120 2.070 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 1.240 0.720 1.640 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 -0.280 2.000 0.280 ;
        RECT  0.800 -0.280 1.880 0.340 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.960 3.320 2.000 3.880 ;
        RECT  0.680 2.560 0.960 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.440 1.360 1.600 1.640 ;
        RECT  1.280 1.290 1.440 2.400 ;
        RECT  1.040 1.290 1.280 1.450 ;
        RECT  0.350 2.240 1.280 2.400 ;
        RECT  0.880 0.910 1.040 1.450 ;
        RECT  0.370 0.910 0.880 1.080 ;
        RECT  0.090 0.800 0.370 1.080 ;
        RECT  0.090 1.940 0.350 2.400 ;
    END
END MAS17

MACRO MAS18
    CLASS CORE ;
    FOREIGN MAS18 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 0.990 2.720 3.000 ;
        RECT  2.430 0.990 2.480 1.270 ;
        RECT  1.650 2.720 2.480 3.000 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.480 0.880 1.750 ;
        RECT  0.480 1.480 0.720 1.960 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.180 1.960 1.620 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 0.440 1.200 0.870 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.070 -0.280 2.800 0.280 ;
        RECT  1.790 -0.280 2.070 0.400 ;
        RECT  0.370 -0.280 1.790 0.280 ;
        RECT  0.090 -0.280 0.370 0.580 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.040 3.320 2.800 3.880 ;
        RECT  1.660 3.200 2.040 3.880 ;
        RECT  0.830 3.260 1.660 3.880 ;
        RECT  0.550 2.680 0.830 3.880 ;
        RECT  0.000 3.320 0.550 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.230 0.480 2.510 0.760 ;
        RECT  1.520 0.600 2.230 0.760 ;
        RECT  2.080 1.970 2.200 2.250 ;
        RECT  1.920 1.970 2.080 2.510 ;
        RECT  1.170 2.350 1.920 2.510 ;
        RECT  1.520 1.910 1.720 2.190 ;
        RECT  1.360 0.600 1.520 2.190 ;
        RECT  0.920 1.030 1.360 1.310 ;
        RECT  0.950 1.970 1.170 2.510 ;
        RECT  0.370 2.350 0.950 2.510 ;
        RECT  0.210 2.350 0.370 2.840 ;
        RECT  0.090 2.560 0.210 2.840 ;
    END
END MAS18

MACRO MAS19
    CLASS CORE ;
    FOREIGN MAS19 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.280 0.440 2.320 1.560 ;
        RECT  2.120 0.440 2.280 2.400 ;
        RECT  2.080 0.440 2.120 1.560 ;
        RECT  2.070 2.080 2.120 2.400 ;
        RECT  2.060 2.120 2.070 2.400 ;
        RECT  1.120 2.120 2.060 2.280 ;
        RECT  0.960 2.120 1.120 2.900 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.640 1.920 1.960 ;
        RECT  1.340 1.640 1.680 1.920 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.520 2.820 2.120 3.000 ;
        RECT  1.280 2.440 1.520 3.000 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.590 0.540 1.900 ;
        RECT  0.340 1.240 0.360 1.900 ;
        RECT  0.080 1.240 0.340 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.880 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.930 -0.280 2.400 0.280 ;
        RECT  0.630 -0.280 0.930 0.760 ;
        RECT  0.000 -0.280 0.630 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.830 3.320 2.400 3.880 ;
        RECT  0.390 3.260 1.830 3.880 ;
        RECT  0.110 2.570 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  0.370 0.920 1.500 1.080 ;
        RECT  0.090 0.600 0.370 1.080 ;
    END
END MAS19

MACRO MAS2
    CLASS CORE ;
    FOREIGN MAS2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.690 0.800 1.240 1.080 ;
        RECT  0.690 2.040 0.920 2.410 ;
        RECT  0.530 0.800 0.690 2.410 ;
        RECT  0.480 2.040 0.530 2.410 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.240 0.370 1.810 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.850 1.240 1.160 1.730 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.370 -0.280 1.600 0.280 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.320 1.600 3.880 ;
        RECT  1.160 2.030 1.440 3.880 ;
        RECT  0.400 3.260 1.160 3.880 ;
        RECT  0.120 2.570 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END MAS2

MACRO MAS20
    CLASS CORE ;
    FOREIGN MAS20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        RECT  2.320 1.240 2.480 1.400 ;
        RECT  1.580 2.200 2.480 2.360 ;
        RECT  2.160 0.980 2.320 1.400 ;
        RECT  1.900 0.980 2.160 1.140 ;
        RECT  1.620 0.860 1.900 1.140 ;
        RECT  1.300 2.200 1.580 3.160 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.070 1.760 2.290 2.040 ;
        RECT  1.560 1.880 2.070 2.040 ;
        RECT  1.300 1.640 1.560 2.040 ;
        RECT  1.020 1.620 1.300 2.040 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.620 0.780 1.960 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.700 -0.280 2.800 0.280 ;
        RECT  2.480 -0.280 2.700 0.990 ;
        RECT  1.060 -0.280 2.480 0.280 ;
        RECT  0.780 -0.280 1.060 1.030 ;
        RECT  0.000 -0.280 0.780 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 3.320 2.800 3.880 ;
        RECT  1.820 2.560 2.100 3.880 ;
        RECT  1.060 3.320 1.820 3.880 ;
        RECT  0.780 2.440 1.060 3.880 ;
        RECT  0.000 3.320 0.780 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.720 1.300 2.000 1.580 ;
        RECT  0.540 1.300 1.720 1.460 ;
        RECT  0.320 1.030 0.540 1.460 ;
        RECT  0.320 2.120 0.540 2.400 ;
        RECT  0.260 1.030 0.320 2.400 ;
        RECT  0.160 1.300 0.260 2.400 ;
    END
END MAS20

MACRO MAS21
    CLASS CORE ;
    FOREIGN MAS21 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.560 0.600 2.720 2.290 ;
        RECT  2.500 0.600 2.560 0.760 ;
        RECT  2.320 2.130 2.560 2.290 ;
        RECT  2.040 0.440 2.500 0.760 ;
        RECT  2.080 2.130 2.320 2.760 ;
        RECT  1.370 2.130 2.080 2.290 ;
        RECT  1.080 2.130 1.370 2.440 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 1.240 1.120 1.740 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.450 1.520 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.960 1.780 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.580 0.380 1.860 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.050 -0.280 2.800 0.280 ;
        RECT  0.750 -0.280 1.050 0.700 ;
        RECT  0.000 -0.280 0.750 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.430 3.190 2.710 3.880 ;
        RECT  1.790 3.320 2.430 3.880 ;
        RECT  0.680 3.030 1.790 3.880 ;
        RECT  0.000 3.320 0.680 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.120 0.920 2.400 1.520 ;
        RECT  0.700 0.920 2.120 1.080 ;
        RECT  0.540 0.920 0.700 2.750 ;
        RECT  0.400 0.920 0.540 1.080 ;
        RECT  0.400 2.590 0.540 2.750 ;
        RECT  0.120 0.800 0.400 1.080 ;
        RECT  0.120 2.590 0.400 2.870 ;
    END
END MAS21

MACRO MAS22
    CLASS CORE ;
    FOREIGN MAS22 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.560 0.650 2.720 2.760 ;
        RECT  2.410 0.650 2.560 0.930 ;
        RECT  2.480 1.640 2.560 2.760 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.600 1.940 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.120 1.580 1.480 1.860 ;
        RECT  0.880 1.240 1.120 1.860 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.410 0.720 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.760 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.210 -0.280 2.800 0.280 ;
        RECT  1.930 -0.280 2.210 0.930 ;
        RECT  0.000 -0.280 1.930 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.170 3.320 2.800 3.880 ;
        RECT  1.890 2.520 2.170 3.880 ;
        RECT  1.220 3.320 1.890 3.880 ;
        RECT  0.480 2.840 1.220 3.880 ;
        RECT  0.000 3.320 0.480 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.260 1.160 2.400 1.440 ;
        RECT  2.100 1.160 2.260 2.280 ;
        RECT  1.770 1.160 2.100 1.320 ;
        RECT  1.680 2.120 2.100 2.280 ;
        RECT  1.610 0.920 1.770 1.320 ;
        RECT  1.400 2.120 1.680 2.800 ;
        RECT  0.780 0.920 1.610 1.080 ;
        RECT  0.750 2.120 1.400 2.280 ;
        RECT  0.330 0.800 0.780 1.080 ;
        RECT  0.530 2.120 0.750 2.400 ;
    END
END MAS22

MACRO MAS23
    CLASS CORE ;
    FOREIGN MAS23 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 0.500 2.320 3.160 ;
        RECT  2.000 0.500 2.160 1.310 ;
        RECT  2.080 1.640 2.160 3.160 ;
        RECT  2.000 1.910 2.080 3.160 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.480 1.520 1.960 ;
        RECT  1.280 1.640 1.300 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.580 1.120 2.410 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 1.580 0.720 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 -0.280 2.400 0.280 ;
        RECT  1.480 -0.280 1.760 0.800 ;
        RECT  0.000 -0.280 1.480 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 3.320 2.400 3.880 ;
        RECT  1.480 3.260 1.760 3.880 ;
        RECT  0.890 3.320 1.480 3.880 ;
        RECT  0.580 3.040 0.890 3.880 ;
        RECT  0.000 3.320 0.580 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.840 1.470 1.920 1.750 ;
        RECT  1.680 1.130 1.840 2.880 ;
        RECT  0.520 1.130 1.680 1.290 ;
        RECT  1.340 2.720 1.680 2.880 ;
        RECT  1.060 2.720 1.340 3.000 ;
        RECT  0.550 2.720 1.060 2.880 ;
        RECT  0.390 2.190 0.550 2.880 ;
        RECT  0.240 1.010 0.520 1.290 ;
        RECT  0.200 2.190 0.390 2.350 ;
    END
END MAS23

MACRO MAS24
    CLASS CORE ;
    FOREIGN MAS24 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 0.870 2.320 1.560 ;
        RECT  2.080 0.870 2.240 2.280 ;
        RECT  2.010 0.870 2.080 1.150 ;
        RECT  1.460 2.120 2.080 2.280 ;
        RECT  1.300 2.120 1.460 2.890 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.620 1.380 1.920 1.960 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.360 1.000 1.580 ;
        RECT  0.480 1.360 0.720 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.250 1.620 1.410 1.900 ;
        RECT  1.120 1.740 1.250 1.900 ;
        RECT  0.880 1.740 1.120 2.360 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.430 3.320 2.800 3.880 ;
        RECT  2.150 2.660 2.430 3.880 ;
        RECT  0.430 3.320 2.150 3.880 ;
        RECT  0.120 2.240 0.430 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.490 0.550 2.650 0.990 ;
        RECT  1.690 0.550 2.490 0.710 ;
        RECT  1.530 0.550 1.690 0.990 ;
        RECT  0.770 0.830 1.530 0.990 ;
        RECT  0.610 0.710 0.770 0.990 ;
    END
END MAS24

MACRO MAS25
    CLASS CORE ;
    FOREIGN MAS25 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.930 0.940 2.090 2.850 ;
        RECT  1.890 0.940 1.930 1.100 ;
        RECT  1.680 2.600 1.930 3.160 ;
        RECT  1.610 0.820 1.890 1.100 ;
        RECT  1.590 2.600 1.680 2.880 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.900 1.070 2.120 ;
        RECT  0.480 1.640 0.760 2.120 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 2.840 1.160 3.160 ;
        RECT  0.500 3.000 0.880 3.160 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.050 -0.280 3.200 0.280 ;
        RECT  2.770 -0.280 3.050 0.400 ;
        RECT  0.930 -0.280 2.770 0.340 ;
        RECT  0.650 -0.280 0.930 1.030 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.010 3.320 3.200 3.880 ;
        RECT  2.730 2.100 3.010 3.880 ;
        RECT  0.340 3.320 2.730 3.880 ;
        RECT  0.710 2.510 0.950 2.680 ;
        RECT  0.520 2.510 0.710 2.770 ;
        RECT  0.340 2.610 0.520 2.770 ;
        RECT  0.160 2.610 0.340 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.850 1.360 2.970 1.640 ;
        RECT  2.690 0.560 2.850 1.640 ;
        RECT  2.210 0.560 2.690 0.720 ;
        RECT  2.250 1.030 2.530 2.880 ;
        RECT  2.050 0.500 2.210 0.720 ;
        RECT  1.450 0.500 2.050 0.660 ;
        RECT  1.610 1.260 1.770 2.440 ;
        RECT  1.450 1.260 1.610 1.420 ;
        RECT  1.390 2.280 1.610 2.440 ;
        RECT  1.290 0.500 1.450 1.420 ;
        RECT  1.230 1.580 1.450 1.900 ;
        RECT  1.170 2.280 1.390 2.590 ;
        RECT  1.130 0.750 1.290 1.030 ;
        RECT  1.080 1.580 1.230 1.740 ;
        RECT  0.920 1.320 1.080 1.740 ;
        RECT  0.370 1.320 0.920 1.480 ;
        RECT  0.320 1.030 0.370 1.480 ;
        RECT  0.160 1.030 0.320 2.450 ;
        RECT  0.090 1.030 0.160 1.310 ;
        RECT  0.100 2.170 0.160 2.450 ;
    END
END MAS25

MACRO MAS26
    CLASS CORE ;
    FOREIGN MAS26 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 0.950 2.320 3.160 ;
        RECT  2.070 0.950 2.160 1.210 ;
        RECT  2.080 2.040 2.160 3.160 ;
        RECT  1.940 2.040 2.080 2.520 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.560 1.560 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.820 2.780 1.160 3.160 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.640 0.760 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.890 -0.280 2.400 0.280 ;
        RECT  1.600 -0.280 1.890 0.550 ;
        RECT  0.840 -0.280 1.600 0.280 ;
        RECT  0.560 -0.280 0.840 0.800 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.740 3.320 2.400 3.880 ;
        RECT  1.460 2.210 1.740 3.880 ;
        RECT  0.000 3.320 1.460 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.880 1.480 2.000 1.780 ;
        RECT  1.720 1.060 1.880 1.780 ;
        RECT  1.300 1.060 1.720 1.240 ;
        RECT  1.080 0.520 1.300 1.240 ;
        RECT  1.020 0.520 1.080 2.280 ;
        RECT  0.920 1.090 1.020 2.280 ;
        RECT  0.120 1.090 0.920 1.250 ;
        RECT  0.580 2.120 0.920 2.280 ;
        RECT  0.300 2.120 0.580 2.400 ;
    END
END MAS26

MACRO MAS27
    CLASS CORE ;
    FOREIGN MAS27 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 0.440 2.490 1.190 ;
        RECT  2.240 1.910 2.360 2.600 ;
        RECT  2.080 0.440 2.240 2.600 ;
        RECT  1.090 2.440 2.080 2.600 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.270 1.120 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.540 1.790 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 1.240 0.720 1.680 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 0.440 3.520 1.750 ;
        RECT  2.970 1.470 3.240 1.750 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.970 -0.280 3.600 0.280 ;
        RECT  0.690 -0.280 0.970 0.640 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.840 3.320 3.600 3.880 ;
        RECT  2.560 2.270 2.840 3.880 ;
        RECT  1.770 3.260 2.560 3.880 ;
        RECT  1.490 3.200 1.770 3.880 ;
        RECT  0.890 3.260 1.490 3.880 ;
        RECT  0.610 2.440 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  3.170 1.910 3.450 2.190 ;
        RECT  2.810 1.910 3.170 2.070 ;
        RECT  2.810 1.030 2.950 1.310 ;
        RECT  2.650 1.030 2.810 2.070 ;
        RECT  2.400 1.430 2.650 1.710 ;
        RECT  1.700 0.920 1.920 2.280 ;
        RECT  0.410 0.920 1.700 1.080 ;
        RECT  0.090 2.120 1.700 2.280 ;
        RECT  0.130 0.800 0.410 1.080 ;
    END
END MAS27

MACRO MAS28
    CLASS CORE ;
    FOREIGN MAS28 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.310 1.240 2.320 2.880 ;
        RECT  2.160 1.030 2.310 2.880 ;
        RECT  2.030 1.030 2.160 2.360 ;
        RECT  1.900 2.720 2.160 2.880 ;
        RECT  1.610 2.720 1.900 3.000 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.200 1.520 1.640 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.370 1.240 0.760 1.640 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 2.350 1.180 2.760 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.780 -0.280 2.400 0.280 ;
        RECT  1.500 -0.280 1.780 0.360 ;
        RECT  0.370 -0.280 1.500 0.340 ;
        RECT  0.090 -0.280 0.370 1.080 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.910 3.320 2.400 3.880 ;
        RECT  1.580 3.200 1.910 3.880 ;
        RECT  0.720 3.320 1.580 3.880 ;
        RECT  0.450 2.560 0.720 3.880 ;
        RECT  0.000 3.320 0.450 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.840 0.520 2.110 0.800 ;
        RECT  1.680 0.520 1.840 2.190 ;
        RECT  1.630 0.520 1.680 1.030 ;
        RECT  0.980 0.810 1.630 1.030 ;
        RECT  0.100 1.910 1.380 2.190 ;
    END
END MAS28

MACRO MAS29
    CLASS CORE ;
    FOREIGN MAS29 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 0.920 2.320 2.760 ;
        RECT  2.160 0.800 2.240 2.930 ;
        RECT  1.960 0.800 2.160 1.080 ;
        RECT  2.080 1.640 2.160 2.930 ;
        RECT  1.960 1.910 2.080 2.930 ;
        RECT  1.300 0.920 1.960 1.080 ;
        RECT  1.020 0.800 1.300 1.080 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.320 1.490 1.520 2.360 ;
        RECT  1.280 2.040 1.320 2.360 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.920 1.750 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.240 0.640 1.770 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.330 1.120 2.360 ;
        RECT  0.480 1.980 0.880 2.360 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.720 -0.280 2.400 0.280 ;
        RECT  1.440 -0.280 1.720 0.400 ;
        RECT  0.500 -0.280 1.440 0.340 ;
        RECT  0.220 -0.280 0.500 1.030 ;
        RECT  0.000 -0.280 0.220 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.920 3.320 2.400 3.880 ;
        RECT  0.640 3.200 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.160 2.650 1.440 2.930 ;
        RECT  0.370 2.650 1.160 2.890 ;
        RECT  0.090 2.590 0.370 2.890 ;
    END
END MAS29

MACRO MAS3
    CLASS CORE ;
    FOREIGN MAS3 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.840 2.120 2.120 2.400 ;
        RECT  1.640 0.800 1.920 1.080 ;
        RECT  0.680 2.120 1.840 2.280 ;
        RECT  0.720 0.920 1.640 1.080 ;
        RECT  0.680 0.440 0.720 1.080 ;
        RECT  0.520 0.440 0.680 2.280 ;
        RECT  0.480 0.440 0.520 1.210 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.240 1.120 1.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.380 1.240 1.920 1.560 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.840 2.320 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.600 3.320 2.400 3.880 ;
        RECT  0.320 2.800 0.600 3.880 ;
        RECT  0.000 3.320 0.320 3.880 ;
        END
    END VDD
END MAS3

MACRO MAS30
    CLASS CORE ;
    FOREIGN MAS30 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 0.440 2.320 2.760 ;
        RECT  1.940 0.440 2.160 0.720 ;
        RECT  2.080 1.640 2.160 2.760 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.470 1.420 1.750 ;
        RECT  1.120 0.840 1.280 1.750 ;
        RECT  0.880 0.840 1.120 1.160 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.400 0.910 1.650 ;
        RECT  0.480 1.240 0.720 1.650 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 -0.280 2.400 0.280 ;
        RECT  1.380 -0.280 1.660 0.610 ;
        RECT  0.650 -0.280 1.380 0.280 ;
        RECT  0.370 -0.280 0.650 1.080 ;
        RECT  0.000 -0.280 0.370 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.790 3.320 2.400 3.880 ;
        RECT  1.510 2.230 1.790 3.880 ;
        RECT  0.370 3.320 1.510 3.880 ;
        RECT  0.090 2.520 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.820 1.390 1.920 1.710 ;
        RECT  1.810 1.030 1.820 1.710 ;
        RECT  1.650 1.030 1.810 2.070 ;
        RECT  1.440 1.030 1.650 1.310 ;
        RECT  1.160 1.910 1.650 2.070 ;
        RECT  1.000 1.910 1.160 2.300 ;
    END
END MAS30

MACRO MAS31
    CLASS CORE ;
    FOREIGN MAS31 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 1.640 2.320 2.760 ;
        RECT  2.080 0.920 2.240 2.760 ;
        RECT  1.660 0.920 2.080 1.080 ;
        RECT  2.010 2.080 2.080 2.760 ;
        RECT  1.380 0.800 1.660 1.080 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.920 1.700 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.200 0.320 2.360 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.580 1.050 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.440 1.520 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  1.940 -0.280 2.220 0.760 ;
        RECT  0.530 -0.280 1.940 0.340 ;
        RECT  0.250 -0.280 0.530 0.930 ;
        RECT  0.000 -0.280 0.250 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.330 3.320 2.400 3.880 ;
        RECT  1.050 2.440 1.330 3.880 ;
        RECT  0.370 3.260 1.050 3.880 ;
        RECT  0.090 2.560 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.530 2.120 1.810 2.820 ;
        RECT  0.850 2.120 1.530 2.280 ;
        RECT  0.570 2.120 0.850 2.800 ;
    END
END MAS31

MACRO MAS32
    CLASS CORE ;
    FOREIGN MAS32 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.700 0.440 2.720 2.360 ;
        RECT  2.480 0.440 2.700 3.100 ;
        RECT  2.420 0.440 2.480 1.220 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 2.040 2.320 2.360 ;
        RECT  1.720 1.740 1.880 2.360 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.240 1.920 1.560 ;
        RECT  1.380 1.240 1.640 1.520 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.060 1.200 1.220 1.560 ;
        RECT  0.880 1.200 1.060 1.580 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.740 0.860 2.020 ;
        RECT  0.440 1.640 0.720 2.020 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.220 3.320 2.800 3.880 ;
        RECT  1.940 2.650 2.220 3.880 ;
        RECT  0.000 3.320 1.940 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.240 1.420 2.320 1.700 ;
        RECT  2.080 0.880 2.240 1.700 ;
        RECT  1.780 0.880 2.080 1.040 ;
        RECT  1.500 0.760 1.780 1.040 ;
        RECT  0.860 0.880 1.500 1.040 ;
        RECT  0.580 0.760 0.860 1.040 ;
        RECT  0.380 2.180 0.660 3.010 ;
        RECT  0.280 0.880 0.580 1.040 ;
        RECT  0.280 2.180 0.380 2.340 ;
        RECT  0.120 0.880 0.280 2.340 ;
    END
END MAS32

MACRO MAS33
    CLASS CORE ;
    FOREIGN MAS33 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.440 2.320 2.280 ;
        RECT  1.900 0.920 2.080 1.080 ;
        RECT  1.580 2.120 2.080 2.280 ;
        RECT  1.290 2.120 1.580 2.530 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.920 1.800 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.720 0.440 2.000 ;
        RECT  0.080 0.440 0.320 2.000 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.720 1.360 0.920 1.640 ;
        RECT  0.670 1.240 0.720 1.640 ;
        RECT  0.480 1.240 0.670 1.560 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.160 1.410 1.520 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 3.320 2.400 3.880 ;
        RECT  1.780 2.440 2.060 3.880 ;
        RECT  0.460 3.320 1.780 3.880 ;
        RECT  0.190 2.340 0.460 3.880 ;
        RECT  0.000 3.320 0.190 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.480 0.710 1.640 0.990 ;
        RECT  0.720 0.830 1.480 0.990 ;
        RECT  0.560 0.710 0.720 0.990 ;
    END
END MAS33

MACRO MAS34
    CLASS CORE ;
    FOREIGN MAS34 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.680 1.090 3.920 2.360 ;
        RECT  3.270 1.090 3.680 1.250 ;
        RECT  3.430 2.170 3.680 2.360 ;
        RECT  3.150 2.170 3.430 2.960 ;
        RECT  2.990 0.970 3.270 1.250 ;
        RECT  1.720 2.520 3.150 2.680 ;
        RECT  1.440 2.520 1.720 2.800 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.410 2.850 1.960 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.170 1.640 3.520 2.010 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.520 0.590 1.800 ;
        RECT  0.080 1.520 0.320 2.760 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.450 1.160 1.960 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 1.790 2.320 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.410 1.920 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.370 -0.280 4.000 0.280 ;
        RECT  1.090 -0.280 1.370 0.800 ;
        RECT  0.370 -0.280 1.090 0.280 ;
        RECT  0.090 -0.280 0.370 1.190 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.560 3.320 4.000 3.880 ;
        RECT  2.280 2.840 2.560 3.880 ;
        RECT  0.880 3.320 2.280 3.880 ;
        RECT  0.600 2.320 0.880 3.880 ;
        RECT  0.000 3.320 0.600 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  3.470 0.650 3.750 0.930 ;
        RECT  2.790 0.650 3.470 0.810 ;
        RECT  2.510 0.650 2.790 1.120 ;
        RECT  1.830 0.650 2.510 0.810 ;
        RECT  2.030 0.970 2.310 1.250 ;
        RECT  0.850 1.090 2.030 1.250 ;
        RECT  1.550 0.650 1.830 0.930 ;
        RECT  0.570 0.770 0.850 1.250 ;
    END
END MAS34

MACRO MAS35
    CLASS CORE ;
    FOREIGN MAS35 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.200 2.160 3.480 2.890 ;
        RECT  2.440 2.160 3.200 2.320 ;
        RECT  2.440 1.240 2.720 1.560 ;
        RECT  2.280 1.080 2.440 2.440 ;
        RECT  1.960 1.080 2.280 1.240 ;
        RECT  2.160 2.120 2.280 2.440 ;
        RECT  1.680 0.650 1.960 1.240 ;
        END
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.400 0.640 1.680 ;
        RECT  0.320 1.400 0.360 2.360 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.480 1.120 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.200 1.520 1.680 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 0.440 3.520 1.560 ;
        RECT  3.010 1.200 3.280 1.480 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.640 3.120 2.000 ;
        RECT  2.600 1.720 2.880 2.000 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.500 2.120 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.120 -0.280 3.600 0.280 ;
        RECT  2.840 -0.280 3.120 0.800 ;
        RECT  0.600 -0.280 2.840 0.340 ;
        RECT  0.320 -0.280 0.600 0.970 ;
        RECT  0.000 -0.280 0.320 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 3.320 3.600 3.880 ;
        RECT  1.120 2.610 1.400 3.880 ;
        RECT  0.440 3.320 1.120 3.880 ;
        RECT  0.160 2.610 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.720 2.610 3.000 2.890 ;
        RECT  1.880 2.730 2.720 2.890 ;
        RECT  1.600 2.160 1.880 2.890 ;
        RECT  0.920 2.160 1.600 2.320 ;
        RECT  0.640 2.160 0.920 2.890 ;
    END
END MAS35

MACRO MAS36
    CLASS CORE ;
    FOREIGN MAS36 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.880 2.320 2.700 ;
        RECT  1.920 0.880 2.080 1.160 ;
        RECT  1.760 2.540 2.080 2.700 ;
        RECT  1.600 2.540 1.760 3.140 ;
        RECT  1.480 2.980 1.600 3.140 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 0.840 1.560 1.580 ;
        RECT  1.240 0.840 1.280 1.160 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 0.440 0.790 0.810 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.060 1.640 1.120 1.960 ;
        RECT  0.820 1.640 1.060 2.060 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.360 -0.280 2.400 0.280 ;
        RECT  1.080 -0.280 1.360 0.400 ;
        RECT  0.000 -0.280 1.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.220 3.320 2.400 3.880 ;
        RECT  1.940 3.200 2.220 3.880 ;
        RECT  1.300 3.320 1.940 3.880 ;
        RECT  1.020 2.800 1.300 3.880 ;
        RECT  0.500 3.260 1.020 3.880 ;
        RECT  0.220 3.200 0.500 3.880 ;
        RECT  0.000 3.320 0.220 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.740 1.640 1.900 2.380 ;
        RECT  0.840 2.220 1.740 2.380 ;
        RECT  0.560 2.220 0.840 2.860 ;
        RECT  0.520 2.220 0.560 2.380 ;
        RECT  0.360 0.970 0.520 2.380 ;
        RECT  0.240 0.970 0.360 1.250 ;
    END
END MAS36

MACRO MAS37
    CLASS CORE ;
    FOREIGN MAS37 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.890 0.810 3.120 2.940 ;
        RECT  2.880 0.810 2.890 1.960 ;
        RECT  2.810 2.660 2.890 2.940 ;
        RECT  1.620 2.660 2.810 2.820 ;
        RECT  1.340 2.410 1.620 2.820 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 2.040 2.720 2.500 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.610 0.500 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.730 1.200 1.120 1.560 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 1.600 2.490 1.820 ;
        RECT  2.080 1.600 2.320 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.270 1.640 1.920 2.070 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.200 -0.280 3.200 0.280 ;
        RECT  0.920 -0.280 1.200 0.400 ;
        RECT  0.400 -0.280 0.920 0.280 ;
        RECT  0.120 -0.280 0.400 0.410 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.570 3.320 3.200 3.880 ;
        RECT  2.290 3.200 2.570 3.880 ;
        RECT  0.670 3.260 2.290 3.880 ;
        RECT  0.390 2.250 0.670 3.880 ;
        RECT  0.000 3.320 0.390 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.360 0.920 2.630 1.370 ;
        RECT  1.660 1.200 2.360 1.370 ;
        RECT  1.870 0.640 2.150 1.040 ;
        RECT  0.800 0.640 1.870 0.800 ;
        RECT  1.390 1.020 1.660 1.370 ;
        RECT  0.520 0.640 0.800 0.970 ;
    END
END MAS37

MACRO MAS38
    CLASS CORE ;
    FOREIGN MAS38 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 0.680 2.720 1.960 ;
        RECT  2.470 0.680 2.630 3.160 ;
        RECT  2.250 0.680 2.470 0.940 ;
        RECT  2.270 2.880 2.470 3.160 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.610 2.040 1.920 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.230 1.050 1.520 1.630 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.170 0.430 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.830 2.040 1.120 2.360 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 -0.280 2.800 0.280 ;
        RECT  1.650 -0.280 2.000 0.560 ;
        RECT  0.000 -0.280 1.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.070 3.320 2.800 3.880 ;
        RECT  1.790 2.880 2.070 3.880 ;
        RECT  0.350 3.320 1.790 3.880 ;
        RECT  0.090 2.460 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.140 2.110 2.300 2.720 ;
        RECT  1.170 2.560 2.140 2.720 ;
        RECT  1.970 1.630 2.040 1.870 ;
        RECT  1.810 0.720 1.970 1.870 ;
        RECT  1.370 0.720 1.810 0.880 ;
        RECT  1.760 1.630 1.810 1.870 ;
        RECT  1.090 0.520 1.370 0.880 ;
        RECT  0.890 2.560 1.170 2.840 ;
        RECT  0.370 0.520 1.090 0.680 ;
        RECT  0.670 2.560 0.890 2.720 ;
        RECT  0.670 0.990 0.750 1.880 ;
        RECT  0.590 0.990 0.670 2.720 ;
        RECT  0.510 1.720 0.590 2.720 ;
        RECT  0.090 0.440 0.370 0.680 ;
    END
END MAS38

MACRO MAS39
    CLASS CORE ;
    FOREIGN MAS39 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 1.240 2.320 2.360 ;
        RECT  2.080 0.840 2.240 2.360 ;
        RECT  0.890 0.840 2.080 1.000 ;
        RECT  1.810 2.120 2.080 2.280 ;
        RECT  1.530 2.120 1.810 2.780 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.720 0.590 1.960 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.640 ;
        RECT  0.480 1.240 0.880 1.560 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.920 1.850 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.280 1.520 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 -0.280 2.400 0.280 ;
        RECT  1.800 -0.280 2.080 0.680 ;
        RECT  0.370 -0.280 1.800 0.290 ;
        RECT  0.090 -0.280 0.370 0.970 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.850 3.320 2.400 3.880 ;
        RECT  0.570 3.250 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.170 2.570 2.290 2.850 ;
        RECT  2.010 2.570 2.170 3.100 ;
        RECT  1.330 2.940 2.010 3.100 ;
        RECT  1.170 2.120 1.330 3.100 ;
        RECT  1.050 2.120 1.170 2.850 ;
        RECT  0.640 2.120 1.050 2.280 ;
        RECT  0.480 2.120 0.640 2.680 ;
        RECT  0.370 2.520 0.480 2.680 ;
        RECT  0.090 2.520 0.370 2.850 ;
    END
END MAS39

MACRO MAS4
    CLASS CORE ;
    FOREIGN MAS4 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.360 1.030 3.520 3.160 ;
        RECT  3.200 1.030 3.360 1.310 ;
        RECT  3.200 1.930 3.360 3.160 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.360 0.720 1.960 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.140 1.140 1.560 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.440 1.210 2.720 1.670 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.040 -0.280 3.600 0.280 ;
        RECT  2.760 -0.280 3.040 0.350 ;
        RECT  0.930 -0.280 2.760 0.340 ;
        RECT  0.650 -0.280 0.930 0.940 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.000 3.320 3.600 3.880 ;
        RECT  2.720 2.670 3.000 3.880 ;
        RECT  0.970 3.260 2.720 3.880 ;
        RECT  0.690 2.500 0.970 3.880 ;
        RECT  0.000 3.320 0.690 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  3.040 1.470 3.200 1.750 ;
        RECT  2.880 0.510 3.040 2.470 ;
        RECT  1.960 0.510 2.880 0.670 ;
        RECT  2.280 2.310 2.880 2.470 ;
        RECT  2.280 0.830 2.440 1.050 ;
        RECT  2.280 1.930 2.410 2.150 ;
        RECT  2.120 0.830 2.280 2.150 ;
        RECT  2.120 2.310 2.280 2.520 ;
        RECT  1.930 2.360 2.120 2.520 ;
        RECT  1.760 0.510 1.960 0.950 ;
        RECT  1.800 1.110 1.960 2.200 ;
        RECT  1.650 2.360 1.930 2.640 ;
        RECT  1.520 1.110 1.800 1.270 ;
        RECT  1.450 2.040 1.800 2.200 ;
        RECT  1.680 0.670 1.760 0.950 ;
        RECT  1.360 1.430 1.640 1.880 ;
        RECT  1.360 0.670 1.520 1.270 ;
        RECT  1.290 2.040 1.450 2.720 ;
        RECT  1.170 0.670 1.360 0.950 ;
        RECT  1.080 1.720 1.360 1.880 ;
        RECT  1.170 2.440 1.290 2.720 ;
        RECT  0.920 1.720 1.080 2.280 ;
        RECT  0.320 2.120 0.920 2.280 ;
        RECT  0.160 0.720 0.320 2.280 ;
        RECT  0.090 0.720 0.160 1.070 ;
        RECT  0.100 2.000 0.160 2.280 ;
    END
END MAS4

MACRO MAS40
    CLASS CORE ;
    FOREIGN MAS40 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.270 0.840 2.320 1.160 ;
        RECT  2.110 0.840 2.270 2.620 ;
        RECT  1.350 0.840 2.110 1.160 ;
        RECT  1.950 2.290 2.110 2.620 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.240 2.720 2.360 ;
        RECT  2.430 1.720 2.480 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.670 1.600 1.950 1.980 ;
        END
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.410 0.320 2.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.810 1.720 0.970 2.360 ;
        RECT  0.480 2.040 0.810 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.190 1.400 1.430 1.680 ;
        RECT  1.150 1.240 1.190 1.680 ;
        RECT  0.880 1.240 1.150 1.560 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.510 -0.280 2.800 0.280 ;
        RECT  2.230 -0.280 2.510 0.680 ;
        RECT  0.470 -0.280 2.230 0.340 ;
        RECT  0.190 -0.280 0.470 1.230 ;
        RECT  0.000 -0.280 0.190 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.230 3.320 2.800 3.880 ;
        RECT  0.180 3.260 1.230 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.430 2.590 2.710 2.950 ;
        RECT  1.750 2.790 2.430 2.950 ;
        RECT  1.470 2.160 1.750 2.950 ;
        RECT  0.850 2.780 1.470 2.950 ;
        RECT  0.540 2.610 0.850 2.950 ;
    END
END MAS40

MACRO MAS41
    CLASS CORE ;
    FOREIGN MAS41 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.740 1.240 8.080 1.640 ;
        RECT  7.580 1.240 7.740 3.160 ;
        RECT  6.820 2.940 7.580 3.160 ;
        END
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.580 1.330 1.960 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.580 0.400 1.860 ;
        RECT  0.080 1.580 0.320 2.760 ;
        END
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.080 1.030 10.320 2.450 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.270 1.030 9.350 1.310 ;
        RECT  9.110 1.030 9.270 2.760 ;
        RECT  8.880 2.440 9.110 2.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.710 2.040 1.920 2.360 ;
        RECT  1.550 1.330 1.710 2.360 ;
        RECT  1.370 2.170 1.550 2.360 ;
        RECT  1.090 2.170 1.370 2.450 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  3.680 1.640 4.120 2.040 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  9.910 -0.280 10.400 0.280 ;
        RECT  9.630 -0.280 9.910 0.420 ;
        RECT  8.470 -0.280 9.630 0.280 ;
        RECT  8.180 -0.280 8.470 0.760 ;
        RECT  3.950 -0.280 8.180 0.280 ;
        RECT  3.670 -0.280 3.950 0.390 ;
        RECT  1.610 -0.280 3.670 0.340 ;
        RECT  1.330 -0.280 1.610 0.400 ;
        RECT  0.350 -0.280 1.330 0.280 ;
        RECT  0.350 1.030 0.400 1.310 ;
        RECT  0.080 -0.280 0.350 1.310 ;
        RECT  0.000 -0.280 0.080 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  9.790 3.320 10.400 3.880 ;
        RECT  9.430 3.240 9.790 3.880 ;
        RECT  8.220 3.320 9.430 3.880 ;
        RECT  7.940 2.460 8.220 3.880 ;
        RECT  6.660 3.320 7.940 3.880 ;
        RECT  6.440 2.850 6.660 3.880 ;
        RECT  5.000 3.320 6.440 3.880 ;
        RECT  4.720 2.990 5.000 3.880 ;
        RECT  3.950 3.320 4.720 3.880 ;
        RECT  3.670 2.990 3.950 3.880 ;
        RECT  1.610 3.260 3.670 3.880 ;
        RECT  1.330 3.200 1.610 3.880 ;
        RECT  0.090 3.260 1.330 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  9.670 1.700 9.790 1.980 ;
        RECT  9.510 0.710 9.670 3.080 ;
        RECT  9.140 0.710 9.510 0.870 ;
        RECT  8.850 2.920 9.510 3.080 ;
        RECT  8.860 0.440 9.140 0.870 ;
        RECT  8.870 1.030 8.950 1.730 ;
        RECT  8.710 1.030 8.870 2.190 ;
        RECT  8.570 2.920 8.850 3.160 ;
        RECT  8.650 1.030 8.710 1.310 ;
        RECT  7.900 1.910 8.710 2.190 ;
        RECT  8.490 1.470 8.520 1.750 ;
        RECT  8.330 0.920 8.490 1.750 ;
        RECT  7.420 0.920 8.330 1.080 ;
        RECT  7.580 0.440 7.860 0.760 ;
        RECT  5.080 0.440 7.580 0.600 ;
        RECT  7.260 0.760 7.420 2.780 ;
        RECT  6.720 0.760 7.260 0.920 ;
        RECT  6.940 2.380 7.260 2.780 ;
        RECT  6.880 1.200 7.100 2.220 ;
        RECT  6.720 2.380 6.940 2.540 ;
        RECT  6.680 1.200 6.880 1.360 ;
        RECT  6.440 1.910 6.720 2.540 ;
        RECT  6.280 1.080 6.680 1.360 ;
        RECT  5.540 0.760 6.440 0.920 ;
        RECT  6.120 1.080 6.280 3.160 ;
        RECT  5.700 1.080 6.120 1.300 ;
        RECT  5.560 3.000 6.120 3.160 ;
        RECT  5.740 1.460 5.960 2.590 ;
        RECT  5.540 1.460 5.740 1.620 ;
        RECT  5.280 2.220 5.560 3.160 ;
        RECT  5.380 0.760 5.540 1.620 ;
        RECT  4.600 1.450 5.380 1.610 ;
        RECT  5.110 1.780 5.330 2.060 ;
        RECT  5.160 2.990 5.280 3.160 ;
        RECT  4.950 1.780 5.110 2.830 ;
        RECT  4.920 0.440 5.080 1.290 ;
        RECT  4.510 2.670 4.950 2.830 ;
        RECT  4.800 1.010 4.920 1.290 ;
        RECT  3.190 2.330 4.790 2.490 ;
        RECT  4.440 1.030 4.600 1.610 ;
        RECT  4.440 1.910 4.560 2.130 ;
        RECT  2.750 0.550 4.510 0.830 ;
        RECT  4.230 2.670 4.510 2.890 ;
        RECT  4.280 1.030 4.440 2.130 ;
        RECT  3.830 1.320 4.280 1.480 ;
        RECT  3.430 2.670 4.230 2.830 ;
        RECT  3.550 1.200 3.830 1.480 ;
        RECT  3.150 2.670 3.430 2.900 ;
        RECT  2.910 0.990 3.190 2.490 ;
        RECT  2.750 2.670 3.150 2.830 ;
        RECT  2.590 0.550 2.750 2.830 ;
        RECT  2.270 0.690 2.430 2.780 ;
        RECT  0.730 0.690 2.270 0.850 ;
        RECT  0.730 2.620 2.270 2.780 ;
        RECT  1.890 1.010 2.110 1.500 ;
        RECT  0.990 1.010 1.890 1.170 ;
        RECT  0.720 1.010 0.990 1.310 ;
        RECT  0.720 2.120 0.930 2.400 ;
        RECT  0.510 0.470 0.730 0.850 ;
        RECT  0.480 2.620 0.730 2.990 ;
        RECT  0.560 1.010 0.720 2.400 ;
    END
END MAS41

MACRO MAS42
    CLASS CORE ;
    FOREIGN MAS42 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.360 1.580 4.720 1.960 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.240 2.320 1.640 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.060 1.580 9.220 2.030 ;
        RECT  8.160 1.640 9.060 2.030 ;
        RECT  7.460 1.870 8.160 2.030 ;
        RECT  7.300 1.380 7.460 2.030 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.520 0.840 11.760 2.650 ;
        RECT  11.280 0.840 11.520 1.960 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  11.270 -0.280 12.000 0.280 ;
        RECT  10.920 -0.280 11.270 0.670 ;
        RECT  9.970 -0.280 10.920 0.280 ;
        RECT  9.690 -0.280 9.970 0.340 ;
        RECT  7.250 -0.280 9.690 0.280 ;
        RECT  6.970 -0.280 7.250 0.340 ;
        RECT  5.730 -0.280 6.970 0.280 ;
        RECT  5.450 -0.280 5.730 0.290 ;
        RECT  4.700 -0.280 5.450 0.280 ;
        RECT  4.420 -0.280 4.700 0.290 ;
        RECT  2.480 -0.280 4.420 0.280 ;
        RECT  2.200 -0.280 2.480 0.290 ;
        RECT  0.840 -0.280 2.200 0.280 ;
        RECT  0.560 -0.280 0.840 0.290 ;
        RECT  0.000 -0.280 0.560 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 3.320 12.000 3.880 ;
        RECT  11.060 2.320 11.300 3.880 ;
        RECT  9.600 3.320 11.060 3.880 ;
        RECT  9.320 2.930 9.600 3.880 ;
        RECT  8.120 3.320 9.320 3.880 ;
        RECT  7.840 3.260 8.120 3.880 ;
        RECT  7.320 3.320 7.840 3.880 ;
        RECT  7.040 3.260 7.320 3.880 ;
        RECT  5.550 3.320 7.040 3.880 ;
        RECT  5.270 3.260 5.550 3.880 ;
        RECT  4.460 3.320 5.270 3.880 ;
        RECT  4.180 3.260 4.460 3.880 ;
        RECT  2.200 3.320 4.180 3.880 ;
        RECT  2.040 2.760 2.200 3.880 ;
        RECT  0.840 3.320 2.040 3.880 ;
        RECT  0.560 3.260 0.840 3.880 ;
        RECT  0.000 3.320 0.560 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  10.900 1.580 11.030 1.860 ;
        RECT  10.740 1.580 10.900 2.540 ;
        RECT  10.500 2.370 10.740 2.540 ;
        RECT  10.420 1.020 10.580 2.190 ;
        RECT  10.200 2.370 10.500 2.670 ;
        RECT  10.340 1.430 10.420 1.710 ;
        RECT  9.860 2.510 10.200 2.670 ;
        RECT  10.020 0.620 10.180 2.210 ;
        RECT  8.510 0.620 10.020 0.780 ;
        RECT  9.700 0.940 9.860 2.670 ;
        RECT  8.360 0.940 9.700 1.100 ;
        RECT  9.160 2.510 9.700 2.670 ;
        RECT  9.380 1.260 9.540 2.350 ;
        RECT  8.180 1.260 9.380 1.420 ;
        RECT  8.620 2.190 9.380 2.350 ;
        RECT  8.880 2.510 9.160 2.730 ;
        RECT  6.050 2.940 8.810 3.100 ;
        RECT  8.460 2.190 8.620 2.470 ;
        RECT  8.230 0.480 8.510 0.780 ;
        RECT  7.660 2.310 8.460 2.470 ;
        RECT  6.670 0.620 8.230 0.780 ;
        RECT  8.020 0.950 8.180 1.420 ;
        RECT  7.940 0.950 8.020 1.230 ;
        RECT  7.780 1.430 7.860 1.710 ;
        RECT  7.620 1.020 7.780 1.710 ;
        RECT  7.500 2.190 7.660 2.470 ;
        RECT  6.990 1.020 7.620 1.180 ;
        RECT  6.960 2.310 7.500 2.470 ;
        RECT  6.960 1.690 7.080 1.980 ;
        RECT  6.830 1.020 6.990 1.250 ;
        RECT  6.800 1.690 6.960 2.470 ;
        RECT  6.430 1.090 6.830 1.250 ;
        RECT  6.510 0.480 6.670 0.930 ;
        RECT  6.040 0.770 6.510 0.930 ;
        RECT  6.210 1.090 6.430 2.370 ;
        RECT  5.720 0.450 6.250 0.610 ;
        RECT  5.890 1.420 6.050 3.100 ;
        RECT  5.880 0.770 6.040 1.250 ;
        RECT  5.550 1.420 5.890 1.580 ;
        RECT  2.520 2.940 5.890 3.100 ;
        RECT  5.040 1.090 5.880 1.250 ;
        RECT  5.570 1.760 5.730 2.040 ;
        RECT  5.560 0.450 5.720 0.930 ;
        RECT  5.100 1.880 5.570 2.040 ;
        RECT  4.200 0.770 5.560 0.930 ;
        RECT  0.640 0.450 5.290 0.610 ;
        RECT  5.040 1.880 5.100 2.690 ;
        RECT  4.880 1.090 5.040 2.690 ;
        RECT  2.840 2.530 4.880 2.690 ;
        RECT  4.040 0.770 4.200 2.360 ;
        RECT  3.690 0.770 4.040 0.930 ;
        RECT  3.420 2.200 4.040 2.360 ;
        RECT  3.660 1.210 3.820 2.040 ;
        RECT  3.530 0.770 3.690 1.050 ;
        RECT  3.360 1.210 3.660 1.370 ;
        RECT  3.600 1.760 3.660 2.040 ;
        RECT  3.200 0.770 3.360 1.370 ;
        RECT  0.960 0.770 3.200 0.930 ;
        RECT  3.040 1.530 3.160 2.370 ;
        RECT  3.000 1.090 3.040 2.370 ;
        RECT  2.880 1.090 3.000 1.690 ;
        RECT  2.740 1.090 2.880 1.310 ;
        RECT  2.680 2.120 2.840 2.690 ;
        RECT  2.120 2.120 2.680 2.280 ;
        RECT  2.360 2.440 2.520 3.100 ;
        RECT  1.800 2.440 2.360 2.600 ;
        RECT  1.960 1.800 2.120 2.280 ;
        RECT  1.600 1.800 1.960 1.960 ;
        RECT  1.640 2.120 1.800 2.600 ;
        RECT  1.460 2.810 1.740 3.090 ;
        RECT  1.280 2.120 1.640 2.280 ;
        RECT  1.440 1.540 1.600 1.960 ;
        RECT  0.960 2.870 1.460 3.030 ;
        RECT  1.280 1.090 1.400 1.310 ;
        RECT  1.120 1.090 1.280 2.280 ;
        RECT  0.800 0.770 0.960 3.030 ;
        RECT  0.480 0.450 0.640 2.830 ;
        RECT  0.120 0.860 0.480 1.080 ;
        RECT  0.090 2.610 0.480 2.830 ;
    END
END MAS42

MACRO MAS43
    CLASS CORE ;
    FOREIGN MAS43 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.060 1.480 7.180 1.640 ;
        RECT  6.900 1.480 7.060 1.930 ;
        RECT  6.240 1.770 6.900 1.930 ;
        RECT  6.120 1.770 6.240 1.980 ;
        RECT  5.960 1.770 6.120 2.360 ;
        RECT  5.520 2.180 5.960 2.360 ;
        RECT  5.420 2.040 5.520 2.360 ;
        RECT  5.260 1.480 5.420 2.360 ;
        RECT  5.120 1.480 5.260 1.640 ;
        END
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.800 2.040 9.920 3.160 ;
        RECT  9.640 0.440 9.800 3.160 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.330 1.240 2.730 1.560 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  0.390 1.240 0.720 1.750 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  9.390 -0.280 10.000 0.280 ;
        RECT  9.100 -0.280 9.390 0.670 ;
        RECT  7.760 -0.280 9.100 0.280 ;
        RECT  7.480 -0.280 7.760 0.340 ;
        RECT  5.160 -0.280 7.480 0.280 ;
        RECT  4.880 -0.280 5.160 0.340 ;
        RECT  3.330 -0.280 4.880 0.280 ;
        RECT  2.530 -0.280 3.330 0.340 ;
        RECT  2.370 -0.280 2.530 1.080 ;
        RECT  0.000 -0.280 2.370 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  9.320 3.320 10.000 3.880 ;
        RECT  9.160 2.930 9.320 3.880 ;
        RECT  7.820 3.320 9.160 3.880 ;
        RECT  7.540 2.850 7.820 3.880 ;
        RECT  6.000 3.320 7.540 3.880 ;
        RECT  5.720 3.260 6.000 3.880 ;
        RECT  5.080 3.320 5.720 3.880 ;
        RECT  4.800 3.260 5.080 3.880 ;
        RECT  2.750 3.320 4.800 3.880 ;
        RECT  2.470 3.260 2.750 3.880 ;
        RECT  0.790 3.320 2.470 3.880 ;
        RECT  0.460 2.660 0.790 3.880 ;
        RECT  0.000 3.320 0.460 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  9.040 1.540 9.200 2.690 ;
        RECT  8.600 2.530 9.040 2.690 ;
        RECT  8.720 0.990 8.880 2.190 ;
        RECT  8.300 0.990 8.720 1.320 ;
        RECT  8.440 2.530 8.600 2.890 ;
        RECT  7.820 2.530 8.440 2.690 ;
        RECT  8.240 1.480 8.400 2.370 ;
        RECT  8.140 1.480 8.240 1.640 ;
        RECT  7.980 0.510 8.140 1.640 ;
        RECT  6.280 0.510 7.980 0.670 ;
        RECT  7.660 0.830 7.820 2.690 ;
        RECT  6.420 0.830 7.660 0.990 ;
        RECT  6.940 2.530 7.660 2.690 ;
        RECT  7.340 1.160 7.500 2.370 ;
        RECT  6.740 1.160 7.340 1.320 ;
        RECT  7.260 2.090 7.340 2.370 ;
        RECT  6.560 2.090 7.260 2.250 ;
        RECT  6.780 2.410 6.940 2.690 ;
        RECT  6.580 1.160 6.740 1.430 ;
        RECT  3.810 2.940 6.720 3.100 ;
        RECT  6.060 1.270 6.580 1.430 ;
        RECT  6.400 2.090 6.560 2.720 ;
        RECT  6.260 0.830 6.420 1.110 ;
        RECT  6.300 2.210 6.400 2.720 ;
        RECT  4.940 2.560 6.300 2.720 ;
        RECT  6.000 0.440 6.280 0.670 ;
        RECT  5.900 0.840 6.060 1.430 ;
        RECT  5.480 0.510 6.000 0.670 ;
        RECT  5.720 0.840 5.900 1.000 ;
        RECT  5.580 1.160 5.740 1.700 ;
        RECT  4.290 1.160 5.580 1.320 ;
        RECT  5.320 0.510 5.480 0.920 ;
        RECT  4.680 0.760 5.320 0.920 ;
        RECT  4.780 1.760 4.940 2.720 ;
        RECT  4.520 0.500 4.680 0.920 ;
        RECT  3.970 0.760 4.520 0.920 ;
        RECT  4.130 1.160 4.290 2.470 ;
        RECT  3.650 0.440 4.210 0.600 ;
        RECT  3.810 0.760 3.970 0.980 ;
        RECT  3.370 0.820 3.810 0.980 ;
        RECT  3.650 1.560 3.810 3.100 ;
        RECT  3.490 0.440 3.650 0.660 ;
        RECT  3.530 1.560 3.650 1.720 ;
        RECT  1.710 2.940 3.650 3.100 ;
        RECT  3.050 0.500 3.490 0.660 ;
        RECT  3.210 0.820 3.370 2.650 ;
        RECT  2.170 2.490 3.210 2.650 ;
        RECT  2.890 0.500 3.050 2.330 ;
        RECT  2.050 0.460 2.210 0.740 ;
        RECT  2.050 1.590 2.170 2.650 ;
        RECT  1.040 0.580 2.050 0.740 ;
        RECT  2.010 0.950 2.050 2.650 ;
        RECT  1.890 0.950 2.010 1.750 ;
        RECT  1.530 1.470 1.890 1.750 ;
        RECT  1.550 1.910 1.710 3.100 ;
        RECT  1.370 1.910 1.550 2.070 ;
        RECT  1.210 0.920 1.370 2.070 ;
        RECT  0.880 0.580 1.040 2.070 ;
        RECT  0.170 0.920 0.880 1.080 ;
        RECT  0.430 1.910 0.880 2.070 ;
        RECT  0.270 1.910 0.430 2.190 ;
    END
END MAS43

MACRO MAS44
    CLASS CORE ;
    FOREIGN MAS44 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 2.840 2.160 3.160 ;
        END
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.190 1.640 1.470 1.960 ;
        RECT  0.760 1.800 1.190 1.960 ;
        RECT  0.400 1.640 0.760 1.960 ;
        END
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.430 1.360 8.690 1.640 ;
        RECT  8.050 1.360 8.430 1.520 ;
        RECT  7.890 0.470 8.050 1.520 ;
        RECT  6.790 0.470 7.890 0.630 ;
        RECT  6.630 0.470 6.790 1.010 ;
        RECT  6.490 0.850 6.630 1.010 ;
        RECT  6.210 0.850 6.490 1.510 ;
        RECT  6.150 0.850 6.210 1.010 ;
        RECT  5.990 0.440 6.150 1.010 ;
        RECT  4.150 0.440 5.990 0.600 ;
        RECT  3.990 0.440 4.150 0.700 ;
        RECT  2.720 0.540 3.990 0.700 ;
        RECT  2.560 0.540 2.720 1.640 ;
        RECT  2.480 0.840 2.560 1.640 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.270 1.640 10.320 2.390 ;
        RECT  10.110 1.030 10.270 2.390 ;
        RECT  9.870 1.030 10.110 1.310 ;
        RECT  10.080 1.640 10.110 2.390 ;
        RECT  9.870 2.110 10.080 2.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.880 0.840 11.120 3.010 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 2.770 1.200 3.160 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.240 3.290 1.620 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  10.630 -0.280 11.200 0.280 ;
        RECT  10.350 -0.280 10.630 0.860 ;
        RECT  8.490 -0.280 10.350 0.280 ;
        RECT  8.210 -0.280 8.490 0.740 ;
        RECT  6.470 -0.280 8.210 0.280 ;
        RECT  6.310 -0.280 6.470 0.690 ;
        RECT  3.830 -0.280 6.310 0.280 ;
        RECT  2.930 -0.280 3.830 0.340 ;
        RECT  2.650 -0.280 2.930 0.380 ;
        RECT  0.370 -0.280 2.650 0.340 ;
        RECT  0.090 -0.280 0.370 0.800 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  10.630 3.320 11.200 3.880 ;
        RECT  10.350 2.990 10.630 3.880 ;
        RECT  9.270 3.320 10.350 3.880 ;
        RECT  8.990 3.260 9.270 3.880 ;
        RECT  8.170 3.320 8.990 3.880 ;
        RECT  7.890 2.800 8.170 3.880 ;
        RECT  5.670 3.320 7.890 3.880 ;
        RECT  5.390 2.450 5.670 3.880 ;
        RECT  3.630 3.320 5.390 3.880 ;
        RECT  3.350 3.200 3.630 3.880 ;
        RECT  2.600 3.260 3.350 3.880 ;
        RECT  2.320 2.740 2.600 3.880 ;
        RECT  0.720 3.320 2.320 3.880 ;
        RECT  0.440 2.800 0.720 3.880 ;
        RECT  0.000 3.320 0.440 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  10.560 1.530 10.720 2.830 ;
        RECT  9.480 2.670 10.560 2.830 ;
        RECT  9.670 0.450 9.810 0.670 ;
        RECT  9.670 1.670 9.730 1.950 ;
        RECT  9.650 2.230 9.690 2.510 ;
        RECT  9.650 0.450 9.670 1.950 ;
        RECT  9.510 0.450 9.650 2.510 ;
        RECT  9.490 1.410 9.510 2.510 ;
        RECT  9.410 2.230 9.490 2.510 ;
        RECT  9.230 2.670 9.480 2.890 ;
        RECT  9.230 1.030 9.350 1.250 ;
        RECT  9.070 1.030 9.230 3.100 ;
        RECT  8.290 1.900 9.070 2.060 ;
        RECT  8.470 2.940 9.070 3.100 ;
        RECT  8.660 2.220 8.880 2.780 ;
        RECT  7.730 2.220 8.660 2.380 ;
        RECT  8.010 1.780 8.290 2.060 ;
        RECT  7.570 0.790 7.730 2.880 ;
        RECT  7.450 0.790 7.570 1.070 ;
        RECT  7.190 2.720 7.570 2.880 ;
        RECT  7.130 2.310 7.410 2.560 ;
        RECT  6.910 2.720 7.190 2.990 ;
        RECT  6.950 0.790 7.170 1.830 ;
        RECT  6.750 2.310 7.130 2.470 ;
        RECT  6.370 1.670 6.950 1.830 ;
        RECT  6.590 2.310 6.750 2.940 ;
        RECT  5.990 2.780 6.590 2.940 ;
        RECT  6.370 2.340 6.430 2.620 ;
        RECT  6.150 1.670 6.370 2.620 ;
        RECT  5.830 1.170 5.990 2.940 ;
        RECT  5.670 0.760 5.830 1.330 ;
        RECT  4.470 0.760 5.670 0.920 ;
        RECT  5.510 2.010 5.670 2.290 ;
        RECT  5.230 2.010 5.510 2.170 ;
        RECT  5.290 1.080 5.470 1.360 ;
        RECT  5.230 1.080 5.290 1.620 ;
        RECT  5.130 1.080 5.230 3.020 ;
        RECT  5.070 1.460 5.130 3.020 ;
        RECT  4.710 2.860 5.070 3.020 ;
        RECT  4.850 1.080 4.970 1.300 ;
        RECT  4.690 1.080 4.850 2.510 ;
        RECT  4.430 2.860 4.710 3.160 ;
        RECT  4.190 2.350 4.690 2.510 ;
        RECT  4.470 1.380 4.530 1.660 ;
        RECT  4.410 0.760 4.470 1.660 ;
        RECT  3.170 2.860 4.430 3.020 ;
        RECT  4.310 0.760 4.410 2.130 ;
        RECT  4.250 0.980 4.310 2.130 ;
        RECT  4.110 0.980 4.250 1.260 ;
        RECT  3.870 1.910 4.250 2.130 ;
        RECT  3.910 2.350 4.190 2.650 ;
        RECT  2.230 2.350 3.910 2.580 ;
        RECT  3.550 0.860 3.710 2.070 ;
        RECT  3.110 0.860 3.550 1.080 ;
        RECT  3.170 1.910 3.550 2.070 ;
        RECT  2.890 1.910 3.170 2.190 ;
        RECT  2.890 2.740 3.170 3.020 ;
        RECT  0.830 0.500 2.400 0.660 ;
        RECT  2.070 0.820 2.230 2.580 ;
        RECT  1.430 0.820 2.070 0.980 ;
        RECT  1.430 2.360 2.070 2.580 ;
        RECT  1.630 1.220 1.910 2.160 ;
        RECT  0.830 1.220 1.630 1.380 ;
        RECT  0.550 0.500 0.830 0.800 ;
        RECT  0.550 1.030 0.830 1.380 ;
        RECT  0.240 1.220 0.550 1.380 ;
        RECT  0.240 2.120 0.370 2.400 ;
        RECT  0.080 1.220 0.240 2.400 ;
    END
END MAS44

MACRO MAS45
    CLASS CORE ;
    FOREIGN MAS45 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.680 1.240 5.920 1.640 ;
        RECT  5.520 1.240 5.680 3.160 ;
        RECT  4.760 2.940 5.520 3.160 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.080 0.610 8.320 3.140 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.110 1.030 7.270 2.760 ;
        RECT  7.050 1.030 7.110 1.310 ;
        RECT  6.880 2.440 7.110 2.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.370 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.640 2.060 1.960 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.370 -0.280 8.400 0.280 ;
        RECT  6.090 -0.280 6.370 0.680 ;
        RECT  1.890 -0.280 6.090 0.280 ;
        RECT  1.610 -0.280 1.890 0.330 ;
        RECT  0.370 -0.280 1.610 0.280 ;
        RECT  0.090 -0.280 0.370 0.330 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.790 3.320 8.400 3.880 ;
        RECT  7.510 3.260 7.790 3.880 ;
        RECT  6.170 3.320 7.510 3.880 ;
        RECT  5.890 2.460 6.170 3.880 ;
        RECT  4.600 3.320 5.890 3.880 ;
        RECT  4.380 2.850 4.600 3.880 ;
        RECT  2.940 3.320 4.380 3.880 ;
        RECT  2.660 2.990 2.940 3.880 ;
        RECT  1.890 3.320 2.660 3.880 ;
        RECT  1.610 2.990 1.890 3.880 ;
        RECT  0.360 3.260 1.610 3.880 ;
        RECT  0.090 2.770 0.360 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  7.800 1.470 7.920 1.750 ;
        RECT  7.640 0.650 7.800 3.080 ;
        RECT  6.930 0.650 7.640 0.810 ;
        RECT  6.870 2.920 7.640 3.080 ;
        RECT  6.650 0.440 6.930 0.810 ;
        RECT  6.710 0.970 6.890 2.190 ;
        RECT  6.590 2.920 6.870 3.130 ;
        RECT  6.400 0.970 6.710 1.250 ;
        RECT  5.840 1.910 6.710 2.190 ;
        RECT  6.240 1.470 6.490 1.750 ;
        RECT  6.080 0.920 6.240 1.750 ;
        RECT  5.360 0.920 6.080 1.080 ;
        RECT  5.330 0.440 5.610 0.740 ;
        RECT  5.200 0.920 5.360 2.780 ;
        RECT  2.930 0.440 5.330 0.600 ;
        RECT  4.850 0.920 5.200 1.080 ;
        RECT  4.880 2.380 5.200 2.780 ;
        RECT  4.820 1.240 5.040 2.220 ;
        RECT  4.660 2.380 4.880 2.540 ;
        RECT  4.690 0.760 4.850 1.080 ;
        RECT  4.470 1.240 4.820 1.400 ;
        RECT  4.570 0.760 4.690 0.920 ;
        RECT  4.380 1.910 4.660 2.540 ;
        RECT  4.220 1.080 4.470 1.400 ;
        RECT  3.390 0.760 4.290 0.920 ;
        RECT  4.060 1.080 4.220 3.160 ;
        RECT  3.550 1.080 4.060 1.300 ;
        RECT  3.500 3.000 4.060 3.160 ;
        RECT  3.680 1.460 3.900 2.590 ;
        RECT  3.390 1.460 3.680 1.620 ;
        RECT  3.220 2.220 3.500 3.160 ;
        RECT  3.320 0.760 3.390 1.620 ;
        RECT  3.230 0.760 3.320 1.610 ;
        RECT  3.050 1.780 3.270 2.060 ;
        RECT  2.450 1.450 3.230 1.610 ;
        RECT  3.100 2.990 3.220 3.160 ;
        RECT  2.890 1.780 3.050 2.830 ;
        RECT  2.770 0.440 2.930 1.290 ;
        RECT  2.450 2.670 2.890 2.830 ;
        RECT  2.650 1.010 2.770 1.290 ;
        RECT  1.070 2.330 2.730 2.490 ;
        RECT  2.380 1.910 2.500 2.130 ;
        RECT  2.380 1.030 2.450 1.610 ;
        RECT  2.170 2.670 2.450 2.890 ;
        RECT  0.750 0.550 2.410 0.830 ;
        RECT  2.220 1.030 2.380 2.130 ;
        RECT  2.130 1.030 2.220 1.480 ;
        RECT  1.370 2.670 2.170 2.830 ;
        RECT  1.770 1.320 2.130 1.480 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.090 2.670 1.370 2.900 ;
        RECT  0.750 2.670 1.090 2.830 ;
        RECT  0.910 0.990 1.070 2.490 ;
        RECT  0.590 0.550 0.750 2.830 ;
    END
END MAS45

MACRO MAS46
    CLASS CORE ;
    FOREIGN MAS46 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 0.910 2.150 2.760 ;
        RECT  1.650 0.910 1.990 1.190 ;
        RECT  1.640 2.440 1.990 2.760 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.130 1.240 1.160 1.560 ;
        RECT  0.820 1.240 1.130 1.630 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.240 2.440 0.720 2.760 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 -0.280 3.200 0.280 ;
        RECT  2.830 -0.280 3.110 0.400 ;
        RECT  0.970 -0.280 2.830 0.340 ;
        RECT  0.690 -0.280 0.970 1.020 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.070 3.320 3.200 3.880 ;
        RECT  2.790 2.240 3.070 3.880 ;
        RECT  0.930 3.260 2.790 3.880 ;
        RECT  0.650 2.920 0.930 3.880 ;
        RECT  0.000 3.320 0.650 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.910 1.540 3.030 1.820 ;
        RECT  2.750 0.590 2.910 1.820 ;
        RECT  1.490 0.590 2.750 0.750 ;
        RECT  2.310 0.980 2.590 2.950 ;
        RECT  1.670 1.350 1.830 2.270 ;
        RECT  1.490 1.350 1.670 1.510 ;
        RECT  1.450 2.110 1.670 2.270 ;
        RECT  1.290 1.670 1.510 1.950 ;
        RECT  1.330 0.590 1.490 1.510 ;
        RECT  1.170 2.110 1.450 2.590 ;
        RECT  1.170 0.740 1.330 1.020 ;
        RECT  0.450 1.790 1.290 1.950 ;
        RECT  0.410 1.790 0.450 2.280 ;
        RECT  0.250 0.980 0.410 2.280 ;
        RECT  0.090 0.980 0.250 1.260 ;
        RECT  0.130 2.000 0.250 2.280 ;
    END
END MAS46

MACRO MAS47
    CLASS CORE ;
    FOREIGN MAS47 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.840 0.840 1.920 1.960 ;
        RECT  1.680 0.840 1.840 2.560 ;
        RECT  1.370 0.920 1.680 1.080 ;
        RECT  1.530 2.280 1.680 2.560 ;
        RECT  0.970 0.800 1.370 1.080 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.460 1.520 1.960 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.430 0.590 1.740 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.830 1.240 1.120 1.870 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.810 -0.280 2.000 0.280 ;
        RECT  1.530 -0.280 1.810 0.680 ;
        RECT  0.390 -0.280 1.530 0.280 ;
        RECT  0.100 -0.280 0.390 0.680 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.850 3.320 2.000 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.050 2.120 1.330 2.560 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.560 ;
    END
END MAS47

MACRO MAS48
    CLASS CORE ;
    FOREIGN MAS48 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.740 0.910 1.920 2.360 ;
        RECT  1.680 0.910 1.740 2.980 ;
        RECT  0.950 0.910 1.680 1.070 ;
        RECT  1.460 2.040 1.680 2.980 ;
        RECT  0.660 0.910 0.950 1.260 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.540 0.660 1.790 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.520 1.120 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.230 1.520 1.800 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.090 -0.280 1.360 0.550 ;
        RECT  0.410 -0.280 1.090 0.280 ;
        RECT  0.130 -0.280 0.410 0.680 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.590 3.320 2.000 3.880 ;
        RECT  0.300 2.190 0.590 3.880 ;
        RECT  0.000 3.320 0.300 3.880 ;
        END
    END VDD
END MAS48

MACRO MAS49
    CLASS CORE ;
    FOREIGN MAS49 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.150 0.440 2.320 2.720 ;
        RECT  2.080 0.440 2.150 1.560 ;
        RECT  1.090 2.440 2.150 2.720 ;
        RECT  1.850 0.790 2.080 1.070 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.910 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.510 1.590 1.960 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.410 1.550 0.720 1.960 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.970 -0.280 2.400 0.280 ;
        RECT  0.690 -0.280 0.970 1.080 ;
        RECT  0.000 -0.280 0.690 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.780 3.320 2.400 3.880 ;
        RECT  1.480 3.090 1.780 3.880 ;
        RECT  0.890 3.260 1.480 3.880 ;
        RECT  0.610 2.460 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.830 1.760 1.990 2.280 ;
        RECT  0.370 2.120 1.830 2.280 ;
        RECT  0.250 1.030 0.410 1.350 ;
        RECT  0.250 2.120 0.370 2.400 ;
        RECT  0.090 1.030 0.250 2.400 ;
    END
END MAS49

MACRO MAS5
    CLASS CORE ;
    FOREIGN MAS5 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.570 1.920 3.110 ;
        RECT  1.600 0.570 1.760 1.320 ;
        RECT  1.680 1.640 1.760 3.110 ;
        RECT  1.610 2.090 1.680 3.110 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.230 1.120 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.370 1.240 0.720 1.770 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.360 -0.280 2.000 0.280 ;
        RECT  1.080 -0.280 1.360 0.470 ;
        RECT  0.370 -0.280 1.080 0.280 ;
        RECT  0.100 -0.280 0.370 1.040 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.360 3.320 2.000 3.880 ;
        RECT  1.080 2.470 1.360 3.880 ;
        RECT  0.000 3.320 1.080 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.450 1.580 1.520 1.860 ;
        RECT  1.440 1.580 1.450 2.310 ;
        RECT  1.280 0.910 1.440 2.310 ;
        RECT  0.890 0.910 1.280 1.070 ;
        RECT  0.400 2.150 1.280 2.310 ;
        RECT  0.610 0.790 0.890 1.070 ;
        RECT  0.120 1.990 0.400 2.620 ;
    END
END MAS5

MACRO MAS50
    CLASS CORE ;
    FOREIGN MAS50 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.470 6.050 1.520 ;
        RECT  4.810 0.470 5.890 0.630 ;
        RECT  4.650 0.470 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.270 1.640 8.320 2.390 ;
        RECT  8.150 1.150 8.270 2.390 ;
        RECT  8.110 1.030 8.150 2.390 ;
        RECT  7.870 1.030 8.110 1.310 ;
        RECT  8.080 1.640 8.110 2.390 ;
        RECT  7.850 2.110 8.080 2.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.830 0.840 9.120 2.190 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.670 -0.280 9.200 0.280 ;
        RECT  8.390 -0.280 8.670 0.400 ;
        RECT  6.490 -0.280 8.390 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.580 3.320 9.200 3.880 ;
        RECT  7.290 3.200 8.580 3.880 ;
        RECT  6.080 3.320 7.290 3.880 ;
        RECT  5.800 3.200 6.080 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  8.640 2.600 8.920 2.880 ;
        RECT  7.010 2.680 8.640 2.880 ;
        RECT  7.670 1.670 7.730 1.950 ;
        RECT  7.670 0.450 7.710 0.670 ;
        RECT  7.650 0.450 7.670 1.950 ;
        RECT  7.510 0.450 7.650 2.520 ;
        RECT  7.430 0.450 7.510 0.670 ;
        RECT  7.490 1.410 7.510 2.520 ;
        RECT  7.370 2.240 7.490 2.520 ;
        RECT  7.010 1.030 7.350 1.250 ;
        RECT  6.850 1.030 7.010 3.160 ;
        RECT  6.290 1.900 6.850 2.060 ;
        RECT  6.260 2.940 6.850 3.160 ;
        RECT  6.470 2.500 6.690 2.780 ;
        RECT  5.730 2.500 6.470 2.660 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 0.790 5.730 2.880 ;
        RECT  5.450 0.790 5.570 1.070 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.970 0.790 5.190 1.830 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.970 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.660 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END MAS50

MACRO MAS51
    CLASS CORE ;
    FOREIGN MAS51 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.680 1.240 6.080 1.640 ;
        RECT  5.520 1.240 5.680 3.160 ;
        RECT  4.760 2.940 5.520 3.160 ;
        END
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.030 1.030 8.320 2.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.270 1.090 7.330 1.250 ;
        RECT  7.050 1.090 7.270 2.760 ;
        RECT  6.880 2.440 7.050 2.760 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.370 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.610 1.640 2.060 1.980 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.380 -0.280 8.400 0.280 ;
        RECT  6.100 -0.280 6.380 0.700 ;
        RECT  1.890 -0.280 6.100 0.280 ;
        RECT  1.610 -0.280 1.890 0.330 ;
        RECT  0.370 -0.280 1.610 0.280 ;
        RECT  0.090 -0.280 0.370 0.330 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.940 3.320 8.400 3.880 ;
        RECT  7.570 3.260 7.940 3.880 ;
        RECT  6.210 3.320 7.570 3.880 ;
        RECT  5.930 2.800 6.210 3.880 ;
        RECT  4.600 3.320 5.930 3.880 ;
        RECT  4.380 2.850 4.600 3.880 ;
        RECT  2.940 3.320 4.380 3.880 ;
        RECT  2.660 2.990 2.940 3.880 ;
        RECT  1.890 3.320 2.660 3.880 ;
        RECT  1.610 2.990 1.890 3.880 ;
        RECT  0.370 3.260 1.610 3.880 ;
        RECT  0.090 2.770 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  7.690 0.710 7.870 3.080 ;
        RECT  7.080 0.710 7.690 0.870 ;
        RECT  6.870 2.920 7.690 3.080 ;
        RECT  6.800 0.440 7.080 0.870 ;
        RECT  6.710 1.030 6.890 2.190 ;
        RECT  6.590 2.920 6.870 3.130 ;
        RECT  6.590 1.030 6.710 1.310 ;
        RECT  5.840 1.910 6.710 2.190 ;
        RECT  6.430 1.470 6.490 1.750 ;
        RECT  6.270 0.920 6.430 1.750 ;
        RECT  5.360 0.920 6.270 1.080 ;
        RECT  5.520 0.440 5.800 0.760 ;
        RECT  3.020 0.440 5.520 0.600 ;
        RECT  5.200 0.760 5.360 2.780 ;
        RECT  4.660 0.760 5.200 0.920 ;
        RECT  4.880 2.380 5.200 2.780 ;
        RECT  4.820 1.200 5.040 2.220 ;
        RECT  4.660 2.380 4.880 2.540 ;
        RECT  4.620 1.200 4.820 1.360 ;
        RECT  4.380 1.910 4.660 2.540 ;
        RECT  4.220 1.080 4.620 1.360 ;
        RECT  3.480 0.760 4.380 0.920 ;
        RECT  4.060 1.080 4.220 3.160 ;
        RECT  3.640 1.080 4.060 1.300 ;
        RECT  3.500 3.000 4.060 3.160 ;
        RECT  3.680 1.460 3.900 2.590 ;
        RECT  3.480 1.460 3.680 1.620 ;
        RECT  3.220 2.220 3.500 3.160 ;
        RECT  3.320 0.760 3.480 1.620 ;
        RECT  2.540 1.450 3.320 1.610 ;
        RECT  3.050 1.780 3.270 2.060 ;
        RECT  3.100 2.990 3.220 3.160 ;
        RECT  2.890 1.780 3.050 2.830 ;
        RECT  2.860 0.440 3.020 1.290 ;
        RECT  2.450 2.670 2.890 2.830 ;
        RECT  2.740 1.010 2.860 1.290 ;
        RECT  1.070 2.330 2.730 2.490 ;
        RECT  2.380 1.030 2.540 1.610 ;
        RECT  2.380 1.910 2.500 2.130 ;
        RECT  0.750 0.550 2.450 0.830 ;
        RECT  2.170 2.670 2.450 2.890 ;
        RECT  2.220 1.030 2.380 2.130 ;
        RECT  1.770 1.320 2.220 1.480 ;
        RECT  1.370 2.670 2.170 2.830 ;
        RECT  1.490 1.200 1.770 1.480 ;
        RECT  1.090 2.670 1.370 2.900 ;
        RECT  0.750 2.670 1.090 2.830 ;
        RECT  0.910 0.990 1.070 2.490 ;
        RECT  0.590 0.550 0.750 2.830 ;
    END
END MAS51

MACRO MAS52
    CLASS CORE ;
    FOREIGN MAS52 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.840 1.120 2.470 ;
        RECT  0.770 1.070 0.880 1.310 ;
        RECT  0.730 2.170 0.880 2.470 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.350 1.520 0.720 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.490 -0.280 1.200 0.280 ;
        RECT  0.210 -0.280 0.490 1.310 ;
        RECT  0.000 -0.280 0.210 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.520 3.320 1.200 3.880 ;
        RECT  0.210 2.170 0.520 3.880 ;
        RECT  0.000 3.320 0.210 3.880 ;
        END
    END VDD
END MAS52

MACRO MAS53
    CLASS CORE ;
    FOREIGN MAS53 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 1.150 2.320 2.370 ;
        RECT  2.080 1.150 2.240 2.680 ;
        RECT  1.830 1.150 2.080 1.310 ;
        RECT  1.350 2.520 2.080 2.680 ;
        RECT  1.550 1.030 1.830 1.310 ;
        RECT  1.070 2.120 1.350 2.870 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.330 1.560 0.540 1.880 ;
        RECT  0.320 1.240 0.330 1.880 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 1.360 1.020 1.640 ;
        RECT  0.700 1.360 0.860 2.360 ;
        RECT  0.480 2.040 0.700 2.360 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.480 1.920 2.360 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.540 1.520 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.830 -0.280 2.400 0.280 ;
        RECT  0.550 -0.280 0.830 0.400 ;
        RECT  0.000 -0.280 0.550 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.230 3.320 2.400 3.880 ;
        RECT  1.950 2.840 2.230 3.880 ;
        RECT  0.510 3.260 1.950 3.880 ;
        RECT  0.230 2.800 0.510 3.880 ;
        RECT  0.000 3.320 0.230 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.030 0.710 2.310 0.990 ;
        RECT  1.350 0.710 2.030 0.870 ;
        RECT  1.190 0.710 1.350 1.060 ;
        RECT  0.150 0.840 1.190 1.060 ;
    END
END MAS53

MACRO MAS54
    CLASS CORE ;
    FOREIGN MAS54 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.740 1.920 3.160 ;
        RECT  1.480 0.740 1.760 1.020 ;
        RECT  1.680 2.040 1.760 3.160 ;
        RECT  0.590 2.320 1.680 2.540 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.380 0.680 1.660 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.120 1.720 1.160 2.000 ;
        RECT  0.880 1.600 1.120 2.000 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.520 1.470 1.600 1.750 ;
        RECT  1.320 1.240 1.520 1.750 ;
        RECT  1.280 1.240 1.320 1.560 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.640 -0.280 2.000 0.280 ;
        RECT  0.360 -0.280 0.640 0.990 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 3.320 2.000 3.880 ;
        RECT  0.120 3.010 1.410 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
END MAS54

MACRO MAS55
    CLASS CORE ;
    FOREIGN MAS55 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.500 1.920 3.160 ;
        RECT  1.600 0.500 1.760 1.310 ;
        RECT  1.680 1.640 1.760 3.160 ;
        RECT  1.600 1.910 1.680 3.160 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.370 1.380 0.720 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 -0.280 2.000 0.280 ;
        RECT  1.110 -0.280 1.410 0.760 ;
        RECT  0.000 -0.280 1.110 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 3.320 2.000 3.880 ;
        RECT  1.120 2.560 1.400 3.880 ;
        RECT  0.390 3.290 1.120 3.880 ;
        RECT  0.130 2.160 0.390 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.440 1.470 1.520 1.750 ;
        RECT  1.280 0.920 1.440 2.340 ;
        RECT  0.430 0.920 1.280 1.080 ;
        RECT  0.830 2.180 1.280 2.340 ;
        RECT  0.670 2.180 0.830 3.000 ;
        RECT  0.550 2.720 0.670 3.000 ;
        RECT  0.150 0.920 0.430 1.220 ;
    END
END MAS55

MACRO MAS56
    CLASS CORE ;
    FOREIGN MAS56 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 0.920 3.120 2.870 ;
        RECT  1.670 0.920 2.880 1.080 ;
        RECT  0.990 0.800 1.670 1.080 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.240 2.720 1.960 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.240 1.010 1.560 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.240 2.320 1.650 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.810 1.560 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.540 -0.280 3.200 0.280 ;
        RECT  2.260 -0.280 2.540 0.740 ;
        RECT  0.430 -0.280 2.260 0.280 ;
        RECT  0.150 -0.280 0.430 0.550 ;
        RECT  0.000 -0.280 0.150 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.330 3.320 3.200 3.880 ;
        RECT  1.050 2.760 1.330 3.880 ;
        RECT  0.350 3.260 1.050 3.880 ;
        RECT  0.090 2.200 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.350 2.120 2.630 2.740 ;
        RECT  1.610 2.440 2.350 2.600 ;
        RECT  1.990 2.120 2.150 2.280 ;
        RECT  1.830 1.810 1.990 2.280 ;
        RECT  0.850 1.810 1.830 1.970 ;
        RECT  1.450 2.130 1.610 2.600 ;
        RECT  0.570 1.810 0.850 2.820 ;
    END
END MAS56

MACRO MAS57
    CLASS CORE ;
    FOREIGN MAS57 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.120 0.800 3.400 1.080 ;
        RECT  3.120 2.650 3.390 2.930 ;
        RECT  3.060 0.920 3.120 1.080 ;
        RECT  3.060 2.040 3.120 2.930 ;
        RECT  2.880 0.920 3.060 2.930 ;
        RECT  1.620 0.920 2.880 1.080 ;
        RECT  1.310 0.800 1.620 1.080 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.420 1.240 0.720 1.620 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.490 1.120 2.000 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 1.240 2.320 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.880 1.560 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.240 2.720 1.620 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 1.240 3.520 2.360 ;
        RECT  3.260 1.240 3.280 1.500 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.560 -0.280 3.600 0.280 ;
        RECT  2.280 -0.280 2.560 0.760 ;
        RECT  0.740 -0.280 2.280 0.280 ;
        RECT  0.460 -0.280 0.740 1.080 ;
        RECT  0.000 -0.280 0.460 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.230 3.320 3.600 3.880 ;
        RECT  0.920 3.240 1.230 3.880 ;
        RECT  0.370 3.320 0.920 3.880 ;
        RECT  0.090 2.890 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.410 2.770 2.680 3.050 ;
        RECT  0.860 2.160 2.090 2.320 ;
        RECT  0.590 2.160 0.860 2.440 ;
    END
END MAS57

MACRO MAS58
    CLASS CORE ;
    FOREIGN MAS58 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 0.940 2.320 3.160 ;
        RECT  1.820 0.940 2.160 1.100 ;
        RECT  2.070 1.910 2.160 3.160 ;
        RECT  2.000 1.910 2.070 2.770 ;
        RECT  1.540 0.820 1.820 1.100 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.580 1.520 1.960 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.580 1.120 2.360 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.230 1.580 0.720 1.960 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.220 -0.280 2.400 0.280 ;
        RECT  0.420 -0.280 2.220 0.340 ;
        RECT  0.140 -0.280 0.420 0.750 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.820 3.320 2.400 3.880 ;
        RECT  1.360 3.260 1.820 3.880 ;
        RECT  1.060 2.860 1.360 3.880 ;
        RECT  0.370 3.260 1.060 3.880 ;
        RECT  0.000 3.320 0.370 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.840 1.260 2.000 1.610 ;
        RECT  1.680 1.260 1.840 2.680 ;
        RECT  1.040 1.260 1.680 1.420 ;
        RECT  0.500 2.520 1.680 2.680 ;
        RECT  0.880 1.000 1.040 1.420 ;
        RECT  0.580 1.000 0.880 1.280 ;
        RECT  0.220 2.120 0.500 2.680 ;
    END
END MAS58

MACRO MAS59
    CLASS CORE ;
    FOREIGN MAS59 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.650 0.770 6.720 3.010 ;
        RECT  6.560 0.440 6.650 3.010 ;
        RECT  6.490 0.440 6.560 0.930 ;
        RECT  6.480 2.440 6.560 3.010 ;
        RECT  5.610 0.770 6.490 0.930 ;
        RECT  6.080 2.440 6.480 2.760 ;
        RECT  5.450 0.450 5.610 0.930 ;
        RECT  5.150 0.450 5.450 0.610 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  2.040 2.040 2.320 2.360 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.110 -0.280 6.800 0.280 ;
        RECT  5.830 -0.280 6.110 0.610 ;
        RECT  4.060 -0.280 5.830 0.280 ;
        RECT  3.900 -0.280 4.060 0.700 ;
        RECT  2.580 -0.280 3.900 0.280 ;
        RECT  1.860 -0.280 2.580 0.640 ;
        RECT  0.400 -0.280 1.860 0.280 ;
        RECT  0.120 -0.280 0.400 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.220 3.320 6.800 3.880 ;
        RECT  5.940 2.920 6.220 3.880 ;
        RECT  4.140 3.320 5.940 3.880 ;
        RECT  3.850 3.260 4.140 3.880 ;
        RECT  2.920 3.320 3.850 3.880 ;
        RECT  2.640 3.260 2.920 3.880 ;
        RECT  1.940 3.320 2.640 3.880 ;
        RECT  1.660 3.260 1.940 3.880 ;
        RECT  0.400 3.320 1.660 3.880 ;
        RECT  0.120 3.260 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  6.240 1.090 6.400 2.230 ;
        RECT  6.120 1.090 6.240 1.250 ;
        RECT  6.120 1.800 6.240 2.230 ;
        RECT  5.640 1.800 6.120 1.960 ;
        RECT  5.820 1.350 5.980 1.640 ;
        RECT  5.180 1.350 5.820 1.510 ;
        RECT  5.380 1.680 5.640 1.960 ;
        RECT  5.020 1.030 5.180 3.160 ;
        RECT  4.850 1.030 5.020 1.310 ;
        RECT  4.830 0.570 4.990 0.870 ;
        RECT  4.700 1.660 4.860 2.990 ;
        RECT  4.690 0.710 4.830 0.870 ;
        RECT  4.690 1.660 4.700 1.940 ;
        RECT  2.340 2.830 4.700 2.990 ;
        RECT  4.530 0.710 4.690 1.940 ;
        RECT  4.380 2.110 4.540 2.670 ;
        RECT  4.110 1.660 4.530 1.940 ;
        RECT  3.950 2.110 4.380 2.270 ;
        RECT  3.240 2.510 4.380 2.670 ;
        RECT  4.190 1.000 4.350 1.310 ;
        RECT  3.950 1.150 4.190 1.310 ;
        RECT  3.790 1.150 3.950 2.270 ;
        RECT  3.470 0.690 3.630 2.270 ;
        RECT  3.410 0.690 3.470 0.850 ;
        RECT  3.250 0.440 3.410 0.850 ;
        RECT  3.240 1.110 3.310 1.880 ;
        RECT  2.910 0.440 3.250 0.600 ;
        RECT  3.150 1.110 3.240 2.670 ;
        RECT  3.080 1.720 3.150 2.670 ;
        RECT  1.770 1.720 3.080 1.880 ;
        RECT  1.160 1.400 2.990 1.560 ;
        RECT  1.660 1.020 2.470 1.180 ;
        RECT  2.180 2.520 2.340 2.990 ;
        RECT  1.360 2.830 2.180 2.990 ;
        RECT  1.610 1.720 1.770 2.000 ;
        RECT  1.500 0.590 1.660 1.180 ;
        RECT  0.800 0.590 1.500 0.750 ;
        RECT  1.200 2.830 1.360 3.110 ;
        RECT  0.800 2.830 1.200 2.990 ;
        RECT  1.130 1.400 1.160 2.670 ;
        RECT  1.000 0.930 1.130 2.670 ;
        RECT  0.970 0.930 1.000 1.560 ;
        RECT  0.640 0.590 0.800 2.990 ;
    END
END MAS59

MACRO MAS6
    CLASS CORE ;
    FOREIGN MAS6 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.840 1.640 1.920 2.760 ;
        RECT  1.680 1.030 1.840 2.760 ;
        RECT  1.560 1.030 1.680 1.310 ;
        RECT  1.240 2.520 1.680 2.680 ;
        RECT  0.960 2.520 1.240 2.810 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.520 1.520 2.360 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.640 0.600 1.960 ;
        RECT  0.080 1.640 0.380 2.760 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.920 1.640 1.120 1.960 ;
        RECT  0.760 1.600 0.920 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 -0.280 2.000 0.280 ;
        RECT  0.600 -0.280 0.880 0.990 ;
        RECT  0.000 -0.280 0.600 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.800 3.320 2.000 3.880 ;
        RECT  1.520 2.930 1.800 3.880 ;
        RECT  0.400 3.320 1.520 3.880 ;
        RECT  0.130 2.920 0.400 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.080 1.030 1.360 1.310 ;
        RECT  0.400 1.150 1.080 1.310 ;
        RECT  0.120 1.030 0.400 1.310 ;
    END
END MAS6

MACRO MAS60
    CLASS CORE ;
    FOREIGN MAS60 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.610 1.080 8.720 2.450 ;
        RECT  8.450 0.440 8.610 3.130 ;
        RECT  8.330 0.440 8.450 1.240 ;
        RECT  8.330 1.970 8.450 3.130 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.430 0.440 7.590 2.060 ;
        RECT  7.280 1.640 7.430 2.060 ;
        END
    END CO
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.510 2.160 5.920 2.760 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 1.430 0.530 1.720 ;
        RECT  0.320 1.430 0.340 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.440 3.120 2.050 ;
        RECT  2.570 1.440 2.880 1.600 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.130 -0.280 8.800 0.280 ;
        RECT  7.850 -0.280 8.130 1.240 ;
        RECT  6.050 -0.280 7.850 0.280 ;
        RECT  5.770 -0.280 6.050 0.340 ;
        RECT  2.930 -0.280 5.770 0.280 ;
        RECT  2.650 -0.280 2.930 0.600 ;
        RECT  0.890 -0.280 2.650 0.280 ;
        RECT  0.610 -0.280 0.890 0.300 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.130 3.320 8.800 3.880 ;
        RECT  7.850 2.570 8.130 3.880 ;
        RECT  5.910 3.320 7.850 3.880 ;
        RECT  5.630 3.260 5.910 3.880 ;
        RECT  2.930 3.320 5.630 3.880 ;
        RECT  2.650 3.260 2.930 3.880 ;
        RECT  0.890 3.320 2.650 3.880 ;
        RECT  0.610 3.260 0.890 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  8.130 1.530 8.270 1.810 ;
        RECT  7.970 1.530 8.130 2.380 ;
        RECT  7.630 2.220 7.970 2.380 ;
        RECT  7.470 2.220 7.630 2.840 ;
        RECT  6.770 2.680 7.470 2.840 ;
        RECT  6.230 3.000 7.440 3.160 ;
        RECT  7.090 2.360 7.310 2.520 ;
        RECT  7.090 1.020 7.210 1.180 ;
        RECT  6.930 0.500 7.090 2.520 ;
        RECT  5.490 0.500 6.930 0.660 ;
        RECT  6.610 0.900 6.770 2.840 ;
        RECT  6.510 0.900 6.610 1.180 ;
        RECT  6.260 1.330 6.420 2.590 ;
        RECT  6.190 1.330 6.260 1.490 ;
        RECT  6.130 2.300 6.260 2.590 ;
        RECT  6.070 2.940 6.230 3.160 ;
        RECT  6.030 0.820 6.190 1.490 ;
        RECT  5.940 1.650 6.100 1.930 ;
        RECT  5.010 2.940 6.070 3.100 ;
        RECT  5.210 0.820 6.030 0.980 ;
        RECT  5.330 1.650 5.940 1.810 ;
        RECT  5.350 0.440 5.490 0.660 ;
        RECT  5.330 1.140 5.490 1.300 ;
        RECT  3.790 0.440 5.350 0.600 ;
        RECT  5.170 1.140 5.330 2.780 ;
        RECT  5.060 0.760 5.210 0.980 ;
        RECT  4.150 0.760 5.060 0.920 ;
        RECT  4.850 1.140 5.010 3.100 ;
        RECT  4.730 1.140 4.850 2.940 ;
        RECT  4.390 2.780 4.730 2.940 ;
        RECT  4.470 1.200 4.570 2.620 ;
        RECT  4.410 1.080 4.470 2.620 ;
        RECT  4.310 1.080 4.410 1.360 ;
        RECT  4.130 2.460 4.410 2.620 ;
        RECT  4.150 1.700 4.250 1.980 ;
        RECT  3.990 0.760 4.150 2.300 ;
        RECT  3.970 2.460 4.130 3.010 ;
        RECT  3.650 2.140 3.990 2.300 ;
        RECT  2.450 2.850 3.970 3.010 ;
        RECT  3.470 1.700 3.830 1.980 ;
        RECT  3.630 0.440 3.790 1.250 ;
        RECT  3.490 2.140 3.650 2.690 ;
        RECT  2.160 0.760 3.630 0.920 ;
        RECT  2.400 2.530 3.490 2.690 ;
        RECT  3.310 1.090 3.470 1.980 ;
        RECT  2.350 1.090 3.310 1.250 ;
        RECT  2.720 2.210 3.250 2.370 ;
        RECT  2.560 2.030 2.720 2.370 ;
        RECT  2.350 2.030 2.560 2.190 ;
        RECT  2.290 2.850 2.450 3.150 ;
        RECT  2.240 2.350 2.400 2.690 ;
        RECT  2.190 1.090 2.350 2.190 ;
        RECT  1.210 2.990 2.290 3.150 ;
        RECT  2.030 2.350 2.240 2.510 ;
        RECT  2.130 1.090 2.190 1.250 ;
        RECT  2.030 0.710 2.160 0.920 ;
        RECT  1.710 2.670 2.080 2.830 ;
        RECT  1.550 0.710 2.030 0.870 ;
        RECT  1.870 1.390 2.030 2.510 ;
        RECT  1.710 1.030 1.870 1.550 ;
        RECT  1.550 1.710 1.710 2.190 ;
        RECT  1.550 2.510 1.710 2.830 ;
        RECT  1.390 0.710 1.550 1.870 ;
        RECT  1.230 2.510 1.550 2.670 ;
        RECT  1.070 1.030 1.230 2.670 ;
        RECT  1.050 2.940 1.210 3.150 ;
        RECT  0.310 2.940 1.050 3.100 ;
        RECT  0.850 1.360 0.910 1.640 ;
        RECT  0.690 0.460 0.850 2.420 ;
        RECT  0.090 0.460 0.690 0.680 ;
        RECT  0.310 2.260 0.690 2.420 ;
        RECT  0.150 2.260 0.310 3.160 ;
    END
END MAS60

MACRO MAS61
    CLASS CORE ;
    FOREIGN MAS61 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 0.840 1.920 2.420 ;
        RECT  1.600 0.840 1.680 1.130 ;
        RECT  1.600 2.050 1.680 2.420 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.780 1.240 1.120 1.840 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.240 0.610 1.560 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.290 -0.280 2.000 0.280 ;
        RECT  1.020 -0.280 1.290 0.760 ;
        RECT  0.000 -0.280 1.020 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.400 3.320 2.000 3.880 ;
        RECT  1.120 2.320 1.400 3.880 ;
        RECT  0.380 3.320 1.120 3.880 ;
        RECT  0.100 2.120 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.440 1.360 1.520 1.640 ;
        RECT  1.280 0.920 1.440 2.160 ;
        RECT  0.670 0.920 1.280 1.080 ;
        RECT  0.860 2.000 1.280 2.160 ;
        RECT  0.580 2.000 0.860 2.300 ;
        RECT  0.510 0.520 0.670 1.080 ;
        RECT  0.090 0.520 0.510 0.680 ;
    END
END MAS61

MACRO MAS62
    CLASS CORE ;
    FOREIGN MAS62 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.990 0.500 3.120 1.160 ;
        RECT  2.990 1.720 3.050 2.660 ;
        RECT  2.890 0.500 2.990 2.660 ;
        RECT  2.830 0.500 2.890 1.880 ;
        RECT  2.310 2.500 2.890 2.660 ;
        RECT  1.770 0.500 2.830 0.720 ;
        RECT  2.050 2.340 2.310 2.660 ;
        END
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.640 0.440 4.720 1.560 ;
        RECT  4.640 2.060 4.700 2.340 ;
        RECT  4.480 0.440 4.640 2.340 ;
        RECT  4.430 2.060 4.480 2.340 ;
        END
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.660 1.640 3.920 1.960 ;
        RECT  3.370 1.800 3.660 1.960 ;
        RECT  3.210 1.800 3.370 2.980 ;
        RECT  2.070 2.820 3.210 2.980 ;
        RECT  2.150 1.260 2.350 2.180 ;
        RECT  1.890 2.020 2.150 2.180 ;
        RECT  1.890 2.820 2.070 3.100 ;
        RECT  1.730 2.020 1.890 3.100 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 1.190 3.520 1.560 ;
        RECT  3.150 1.340 3.280 1.560 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.140 -0.280 4.800 0.280 ;
        RECT  3.860 -0.280 4.140 0.700 ;
        RECT  3.530 -0.280 3.860 0.280 ;
        RECT  3.250 -0.280 3.530 0.400 ;
        RECT  0.460 -0.280 3.250 0.280 ;
        RECT  0.180 -0.280 0.460 0.340 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.310 3.320 4.800 3.880 ;
        RECT  4.030 3.200 4.310 3.880 ;
        RECT  3.190 3.260 4.030 3.880 ;
        RECT  2.910 3.200 3.190 3.880 ;
        RECT  0.980 3.260 2.910 3.880 ;
        RECT  0.700 3.200 0.980 3.880 ;
        RECT  0.000 3.320 0.700 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  4.240 1.000 4.320 1.560 ;
        RECT  4.080 1.000 4.240 2.280 ;
        RECT  4.070 1.000 4.080 1.160 ;
        RECT  3.750 2.120 4.080 2.280 ;
        RECT  3.790 0.880 4.070 1.160 ;
        RECT  3.530 2.120 3.750 2.400 ;
        RECT  2.670 2.060 2.730 2.340 ;
        RECT  2.510 0.880 2.670 2.340 ;
        RECT  1.990 0.880 2.510 1.100 ;
        RECT  1.830 0.880 1.990 1.860 ;
        RECT  1.010 1.700 1.830 1.860 ;
        RECT  1.450 0.910 1.670 1.540 ;
        RECT  1.290 2.690 1.570 2.990 ;
        RECT  1.240 0.450 1.530 0.730 ;
        RECT  0.630 0.910 1.450 1.190 ;
        RECT  1.140 2.020 1.420 2.530 ;
        RECT  0.310 2.690 1.290 2.850 ;
        RECT  0.310 0.570 1.240 0.730 ;
        RECT  0.630 2.020 1.140 2.180 ;
        RECT  0.790 1.580 1.010 1.860 ;
        RECT  0.470 0.910 0.630 2.180 ;
        RECT  0.090 0.570 0.310 2.850 ;
    END
END MAS62

MACRO MAS63
    CLASS CORE ;
    FOREIGN MAS63 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.330 0.710 3.490 2.760 ;
        RECT  2.210 0.710 3.330 0.870 ;
        RECT  2.480 2.600 3.330 2.760 ;
        RECT  2.040 2.440 2.480 3.110 ;
        RECT  1.930 0.590 2.210 0.870 ;
        RECT  1.290 0.710 1.930 0.870 ;
        RECT  1.010 0.710 1.290 0.990 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.520 1.120 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.160 1.560 1.600 ;
        END
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.760 1.640 3.160 1.960 ;
        END
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.760 -0.280 3.600 0.280 ;
        RECT  2.480 -0.280 2.760 0.400 ;
        RECT  1.690 -0.280 2.480 0.280 ;
        RECT  0.770 -0.280 1.690 0.340 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.170 3.320 3.600 3.880 ;
        RECT  2.890 3.080 3.170 3.880 ;
        RECT  1.040 3.320 2.890 3.880 ;
        RECT  0.760 2.840 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.890 2.120 3.170 2.440 ;
        RECT  2.880 1.030 3.160 1.310 ;
        RECT  2.600 2.120 2.890 2.280 ;
        RECT  2.600 1.140 2.880 1.310 ;
        RECT  2.440 1.140 2.600 2.280 ;
        RECT  2.020 1.140 2.440 1.300 ;
        RECT  2.000 1.580 2.280 1.860 ;
        RECT  1.740 1.140 2.020 1.420 ;
        RECT  1.880 1.700 2.000 1.860 ;
        RECT  1.720 1.700 1.880 2.680 ;
        RECT  0.680 2.490 1.720 2.680 ;
        RECT  0.520 0.920 0.680 2.680 ;
        RECT  0.370 0.920 0.520 1.080 ;
        RECT  0.210 2.520 0.520 2.680 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END MAS63

MACRO MAS64
    CLASS CORE ;
    FOREIGN MAS64 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.310 1.030 3.470 2.940 ;
        RECT  2.760 1.030 3.310 1.190 ;
        RECT  1.890 2.780 3.310 2.940 ;
        RECT  2.480 0.800 2.760 1.190 ;
        RECT  1.970 0.800 2.480 0.960 ;
        RECT  1.690 0.800 1.970 1.080 ;
        RECT  1.610 2.780 1.890 3.060 ;
        RECT  0.850 2.780 1.610 2.940 ;
        RECT  0.570 2.780 0.850 3.060 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.990 1.460 3.150 2.620 ;
        RECT  0.670 2.460 2.990 2.620 ;
        RECT  0.670 1.240 0.720 1.560 ;
        RECT  0.510 1.240 0.670 2.620 ;
        RECT  0.290 1.240 0.510 1.680 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.120 2.140 2.810 2.300 ;
        RECT  0.960 1.640 1.120 2.300 ;
        RECT  0.880 1.640 0.960 1.980 ;
        RECT  0.830 1.720 0.880 1.980 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.560 1.760 2.490 1.920 ;
        RECT  1.280 1.240 1.560 1.920 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.870 1.240 2.320 1.600 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.410 -0.280 3.600 0.280 ;
        RECT  3.130 -0.280 3.410 0.870 ;
        RECT  0.480 -0.280 3.130 0.280 ;
        RECT  0.200 -0.280 0.480 0.990 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.410 3.320 3.600 3.880 ;
        RECT  2.130 3.200 2.410 3.880 ;
        RECT  1.370 3.320 2.130 3.880 ;
        RECT  1.090 3.200 1.370 3.880 ;
        RECT  0.350 3.320 1.090 3.880 ;
        RECT  0.090 2.050 0.350 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
END MAS64

MACRO MAS65
    CLASS CORE ;
    FOREIGN MAS65 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.360 1.440 2.640 3.100 ;
        RECT  1.680 1.440 2.360 2.160 ;
        RECT  1.480 0.890 1.680 3.160 ;
        RECT  1.400 0.890 1.480 1.350 ;
        RECT  1.400 2.060 1.480 3.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.240 0.840 1.560 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.200 -0.280 2.800 0.280 ;
        RECT  1.920 -0.280 2.200 1.080 ;
        RECT  1.160 -0.280 1.920 0.280 ;
        RECT  0.880 -0.280 1.160 0.760 ;
        RECT  0.000 -0.280 0.880 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.160 3.320 2.800 3.880 ;
        RECT  1.880 2.480 2.160 3.880 ;
        RECT  1.200 3.320 1.880 3.880 ;
        RECT  0.920 2.340 1.200 3.880 ;
        RECT  0.000 3.320 0.920 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.160 1.560 1.270 1.840 ;
        RECT  1.000 0.920 1.160 2.070 ;
        RECT  0.640 0.920 1.000 1.080 ;
        RECT  0.720 1.910 1.000 2.070 ;
        RECT  0.440 1.910 0.720 3.040 ;
        RECT  0.360 0.800 0.640 1.080 ;
    END
END MAS65

MACRO MAS66
    CLASS CORE ;
    FOREIGN MAS66 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.800 1.240 1.920 2.360 ;
        RECT  1.640 1.040 1.800 2.360 ;
        RECT  1.440 1.040 1.640 1.200 ;
        RECT  1.430 2.160 1.640 2.360 ;
        RECT  1.160 0.920 1.440 1.200 ;
        RECT  1.130 2.160 1.430 2.870 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.240 0.760 1.640 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.910 -0.280 2.000 0.280 ;
        RECT  1.630 -0.280 1.910 0.870 ;
        RECT  0.930 -0.280 1.630 0.280 ;
        RECT  0.610 -0.280 0.930 1.030 ;
        RECT  0.000 -0.280 0.610 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.600 2.580 1.910 3.880 ;
        RECT  0.910 3.320 1.600 3.880 ;
        RECT  0.610 2.350 0.910 3.880 ;
        RECT  0.000 3.320 0.610 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.270 1.360 1.390 1.680 ;
        RECT  1.100 1.360 1.270 1.960 ;
        RECT  0.380 1.800 1.100 1.960 ;
        RECT  0.260 0.800 0.410 1.080 ;
        RECT  0.260 1.800 0.380 2.690 ;
        RECT  0.100 0.800 0.260 2.690 ;
    END
END MAS66

MACRO MAS67
    CLASS CORE ;
    FOREIGN MAS67 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.430 0.440 10.720 3.160 ;
        END
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 1.450 1.640 1.960 ;
        RECT  1.280 0.540 1.440 1.960 ;
        RECT  0.680 0.540 1.280 0.700 ;
        RECT  0.520 0.470 0.680 0.700 ;
        RECT  0.370 0.470 0.520 0.630 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.240 0.800 1.960 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  3.600 1.040 3.820 1.630 ;
        RECT  3.440 1.470 3.600 1.960 ;
        RECT  3.280 1.640 3.440 1.960 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  10.230 -0.280 10.800 0.280 ;
        RECT  9.950 -0.280 10.230 0.760 ;
        RECT  9.090 -0.280 9.950 0.300 ;
        RECT  3.240 -0.280 9.090 0.280 ;
        RECT  2.960 -0.280 3.240 0.400 ;
        RECT  1.370 -0.280 2.960 0.280 ;
        RECT  1.090 -0.280 1.370 0.380 ;
        RECT  0.000 -0.280 1.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  10.230 3.320 10.800 3.880 ;
        RECT  8.900 2.800 10.230 3.880 ;
        RECT  7.300 3.320 8.900 3.880 ;
        RECT  7.020 3.260 7.300 3.880 ;
        RECT  5.440 3.320 7.020 3.880 ;
        RECT  5.160 3.200 5.440 3.880 ;
        RECT  3.500 3.320 5.160 3.880 ;
        RECT  3.220 3.200 3.500 3.880 ;
        RECT  1.640 3.260 3.220 3.880 ;
        RECT  1.360 3.200 1.640 3.880 ;
        RECT  0.000 3.320 1.360 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  10.070 1.040 10.230 2.050 ;
        RECT  9.640 1.040 10.070 1.200 ;
        RECT  9.640 1.890 10.070 2.050 ;
        RECT  9.630 1.360 9.910 1.640 ;
        RECT  9.360 0.920 9.640 1.200 ;
        RECT  9.360 1.890 9.640 2.210 ;
        RECT  8.830 1.360 9.630 1.520 ;
        RECT  9.150 0.920 9.360 1.080 ;
        RECT  9.210 1.890 9.360 2.050 ;
        RECT  8.990 1.770 9.210 2.050 ;
        RECT  8.990 0.460 9.150 1.080 ;
        RECT  8.340 0.460 8.990 0.620 ;
        RECT  8.670 0.780 8.830 2.460 ;
        RECT  8.180 0.780 8.670 1.000 ;
        RECT  8.020 2.300 8.670 2.460 ;
        RECT  8.230 1.190 8.510 2.130 ;
        RECT  8.230 2.940 8.510 3.160 ;
        RECT  8.180 0.440 8.340 0.620 ;
        RECT  8.020 1.190 8.230 1.410 ;
        RECT  6.750 2.940 8.230 3.100 ;
        RECT  3.680 0.440 8.180 0.600 ;
        RECT  7.860 0.760 8.020 1.410 ;
        RECT  5.240 0.760 7.860 0.920 ;
        RECT  7.700 1.800 7.820 2.720 ;
        RECT  7.540 1.080 7.700 2.720 ;
        RECT  7.400 1.080 7.540 1.240 ;
        RECT  6.910 2.360 7.540 2.640 ;
        RECT  6.960 1.560 7.380 1.720 ;
        RECT  6.800 1.140 6.960 2.190 ;
        RECT  6.120 1.140 6.800 1.320 ;
        RECT  6.120 2.030 6.800 2.190 ;
        RECT  6.590 2.560 6.750 3.100 ;
        RECT  5.960 1.680 6.640 1.840 ;
        RECT  5.960 2.560 6.590 2.720 ;
        RECT  6.210 2.880 6.430 3.160 ;
        RECT  2.520 2.880 6.210 3.040 ;
        RECT  5.800 1.300 5.960 2.720 ;
        RECT  5.680 1.300 5.800 1.460 ;
        RECT  2.840 2.560 5.800 2.720 ;
        RECT  5.400 1.180 5.680 1.460 ;
        RECT  5.240 1.620 5.640 1.900 ;
        RECT  5.080 0.760 5.240 2.280 ;
        RECT  4.610 0.760 5.080 1.060 ;
        RECT  4.300 2.000 5.080 2.280 ;
        RECT  4.140 1.330 4.920 1.610 ;
        RECT  4.140 0.770 4.320 0.990 ;
        RECT  3.980 0.770 4.140 1.970 ;
        RECT  3.760 1.810 3.980 1.970 ;
        RECT  3.520 0.440 3.680 0.720 ;
        RECT  3.440 0.560 3.520 0.720 ;
        RECT  3.280 0.560 3.440 1.310 ;
        RECT  3.000 1.150 3.280 1.430 ;
        RECT  2.900 0.710 3.120 0.990 ;
        RECT  2.840 0.830 2.900 0.990 ;
        RECT  2.680 0.830 2.840 2.720 ;
        RECT  2.360 0.550 2.520 3.040 ;
        RECT  1.680 0.550 2.360 0.830 ;
        RECT  2.240 2.520 2.360 3.040 ;
        RECT  0.420 2.880 2.240 3.040 ;
        RECT  2.080 1.350 2.200 1.630 ;
        RECT  2.080 2.020 2.200 2.300 ;
        RECT  1.920 1.010 2.080 2.720 ;
        RECT  1.600 1.010 1.920 1.290 ;
        RECT  0.680 2.560 1.920 2.720 ;
        RECT  0.960 0.860 1.120 2.400 ;
        RECT  0.570 0.860 0.960 1.080 ;
        RECT  0.840 2.120 0.960 2.400 ;
        RECT  0.520 2.170 0.680 2.720 ;
        RECT  0.400 2.170 0.520 2.450 ;
        RECT  0.360 2.880 0.420 3.140 ;
        RECT  0.240 0.790 0.370 1.070 ;
        RECT  0.240 2.610 0.360 3.140 ;
        RECT  0.080 0.790 0.240 3.140 ;
    END
END MAS67

MACRO MAS68
    CLASS CORE ;
    FOREIGN MAS68 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 1.130 5.120 2.760 ;
        RECT  4.720 1.130 4.880 1.370 ;
        RECT  3.860 2.520 4.880 2.760 ;
        RECT  4.480 0.600 4.720 1.370 ;
        RECT  3.780 0.600 4.480 0.840 ;
        RECT  3.580 2.440 3.860 2.760 ;
        RECT  3.770 0.440 3.780 0.840 ;
        RECT  3.520 0.440 3.770 1.060 ;
        RECT  1.620 2.440 3.580 2.660 ;
        RECT  3.500 0.440 3.520 0.840 ;
        RECT  1.400 0.560 3.500 0.840 ;
        RECT  1.340 2.440 1.620 2.720 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.560 1.720 4.720 2.280 ;
        RECT  4.320 2.120 4.560 2.280 ;
        RECT  4.080 2.040 4.320 2.360 ;
        RECT  2.720 2.120 4.080 2.280 ;
        RECT  2.440 1.720 2.720 2.280 ;
        RECT  0.740 2.120 2.440 2.280 ;
        RECT  0.580 1.680 0.740 2.280 ;
        RECT  0.340 1.680 0.580 1.850 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.160 1.220 4.320 1.700 ;
        RECT  3.480 1.220 4.160 1.400 ;
        RECT  3.360 1.220 3.480 1.640 ;
        RECT  3.200 1.080 3.360 1.640 ;
        RECT  1.960 1.080 3.200 1.240 ;
        RECT  1.680 1.080 1.960 1.640 ;
        RECT  0.890 1.080 1.680 1.240 ;
        RECT  0.600 0.840 0.890 1.460 ;
        RECT  0.480 0.840 0.600 1.160 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.680 1.640 3.920 1.960 ;
        RECT  3.040 1.800 3.680 1.960 ;
        RECT  2.880 1.400 3.040 1.960 ;
        RECT  2.280 1.400 2.880 1.560 ;
        RECT  2.120 1.400 2.280 1.960 ;
        RECT  1.420 1.800 2.120 1.960 ;
        RECT  1.140 1.680 1.420 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.320 -0.280 5.200 0.280 ;
        RECT  4.040 -0.280 4.320 0.400 ;
        RECT  3.260 -0.280 4.040 0.280 ;
        RECT  2.980 -0.280 3.260 0.400 ;
        RECT  2.200 -0.280 2.980 0.280 ;
        RECT  1.920 -0.280 2.200 0.400 ;
        RECT  1.200 -0.280 1.920 0.280 ;
        RECT  0.920 -0.280 1.200 0.670 ;
        RECT  0.000 -0.280 0.920 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  5.020 3.320 5.200 3.880 ;
        RECT  4.740 3.010 5.020 3.880 ;
        RECT  2.740 3.320 4.740 3.880 ;
        RECT  2.460 2.820 2.740 3.880 ;
        RECT  0.420 3.260 2.460 3.880 ;
        RECT  0.140 2.120 0.420 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
END MAS68

MACRO MAS69
    CLASS CORE ;
    FOREIGN MAS69 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.520 0.440 1.810 1.060 ;
        RECT  0.850 0.900 1.520 1.060 ;
        RECT  1.280 2.670 1.520 3.160 ;
        RECT  0.240 2.670 1.280 2.830 ;
        RECT  0.570 0.440 0.850 1.060 ;
        RECT  0.240 0.900 0.570 1.060 ;
        RECT  0.080 0.900 0.240 2.830 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.340 1.580 2.460 1.860 ;
        RECT  2.180 1.580 2.340 2.510 ;
        RECT  0.720 2.350 2.180 2.510 ;
        RECT  0.560 2.040 0.720 2.510 ;
        RECT  0.400 1.840 0.560 2.510 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.810 1.590 1.930 1.750 ;
        RECT  1.650 1.590 1.810 2.180 ;
        RECT  1.040 2.020 1.650 2.180 ;
        RECT  1.040 1.240 1.120 1.580 ;
        RECT  0.880 1.240 1.040 2.180 ;
        RECT  0.690 1.240 0.880 1.580 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 0.440 2.760 0.760 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 -0.280 3.200 0.280 ;
        RECT  2.160 -0.280 2.320 0.820 ;
        RECT  1.330 -0.280 2.160 0.280 ;
        RECT  1.050 -0.280 1.330 0.670 ;
        RECT  0.370 -0.280 1.050 0.280 ;
        RECT  0.090 -0.280 0.370 0.670 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.870 3.320 3.200 3.880 ;
        RECT  2.590 2.920 2.870 3.880 ;
        RECT  0.370 3.320 2.590 3.880 ;
        RECT  0.090 2.990 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.830 0.920 3.110 2.380 ;
        RECT  1.440 1.260 2.830 1.420 ;
        RECT  1.280 1.260 1.440 1.640 ;
    END
END MAS69

MACRO MAS7
    CLASS CORE ;
    FOREIGN MAS7 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.920 0.440 2.140 0.610 ;
        RECT  1.870 0.440 1.920 0.760 ;
        RECT  1.810 0.440 1.870 2.160 ;
        RECT  1.710 0.440 1.810 2.510 ;
        RECT  1.680 0.440 1.710 0.760 ;
        RECT  1.530 2.000 1.710 2.510 ;
        RECT  0.850 2.000 1.530 2.160 ;
        RECT  0.570 2.000 0.850 2.500 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.240 0.590 1.520 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.840 1.120 1.840 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.550 1.840 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.840 2.320 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.680 -0.280 2.400 0.280 ;
        RECT  0.360 -0.280 0.680 0.680 ;
        RECT  0.000 -0.280 0.360 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.280 3.320 2.400 3.880 ;
        RECT  2.000 2.290 2.280 3.880 ;
        RECT  1.320 3.320 2.000 3.880 ;
        RECT  1.040 2.320 1.320 3.880 ;
        RECT  0.360 3.320 1.040 3.880 ;
        RECT  0.080 2.120 0.360 3.880 ;
        RECT  0.000 3.320 0.080 3.880 ;
        END
    END VDD
END MAS7

MACRO MAS70
    CLASS CORE ;
    FOREIGN MAS70 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.080 0.920 8.320 2.420 ;
        RECT  8.000 0.920 8.080 1.200 ;
        RECT  8.000 1.910 8.080 2.420 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.640 0.440 5.960 0.780 ;
        RECT  5.580 0.500 5.640 0.780 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.480 1.580 2.720 1.960 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.200 2.320 1.560 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.240 0.500 1.560 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 1.240 3.580 1.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.360 1.640 5.560 1.960 ;
        RECT  5.240 1.520 5.360 1.960 ;
        RECT  5.140 1.520 5.240 1.800 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.880 -0.280 8.400 0.280 ;
        RECT  7.600 -0.280 7.880 0.400 ;
        RECT  5.420 -0.280 7.600 0.280 ;
        RECT  5.140 -0.280 5.420 0.930 ;
        RECT  3.420 -0.280 5.140 0.340 ;
        RECT  3.200 -0.280 3.420 1.040 ;
        RECT  2.480 -0.280 3.200 0.280 ;
        RECT  2.200 -0.280 2.480 1.040 ;
        RECT  0.460 -0.280 2.200 0.340 ;
        RECT  0.180 -0.280 0.460 0.940 ;
        RECT  0.000 -0.280 0.180 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.880 3.320 8.400 3.880 ;
        RECT  7.600 3.200 7.880 3.880 ;
        RECT  3.380 3.260 7.600 3.880 ;
        RECT  3.100 2.930 3.380 3.880 ;
        RECT  2.540 3.320 3.100 3.880 ;
        RECT  2.260 2.930 2.540 3.880 ;
        RECT  0.460 3.260 2.260 3.880 ;
        RECT  0.180 2.590 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  7.840 1.360 7.920 1.640 ;
        RECT  7.680 0.620 7.840 1.640 ;
        RECT  6.940 0.620 7.680 0.780 ;
        RECT  7.300 0.940 7.420 1.220 ;
        RECT  7.300 2.200 7.420 2.950 ;
        RECT  7.140 0.940 7.300 3.090 ;
        RECT  3.700 2.930 7.140 3.090 ;
        RECT  6.660 0.620 6.940 2.480 ;
        RECT  6.460 1.060 6.500 2.490 ;
        RECT  6.350 0.940 6.460 2.490 ;
        RECT  6.340 0.940 6.350 2.770 ;
        RECT  6.180 0.940 6.340 1.220 ;
        RECT  6.180 2.170 6.340 2.770 ;
        RECT  6.000 1.530 6.180 1.810 ;
        RECT  4.600 2.610 6.180 2.770 ;
        RECT  5.840 0.970 6.000 2.420 ;
        RECT  5.720 0.970 5.840 1.250 ;
        RECT  5.680 2.200 5.840 2.420 ;
        RECT  4.760 0.650 4.980 2.390 ;
        RECT  4.660 0.650 4.760 0.930 ;
        RECT  4.440 1.090 4.600 2.770 ;
        RECT  4.380 1.090 4.440 1.250 ;
        RECT  4.100 2.610 4.440 2.770 ;
        RECT  4.100 0.910 4.380 1.250 ;
        RECT  4.120 1.410 4.280 2.450 ;
        RECT  3.900 1.410 4.120 1.570 ;
        RECT  3.620 2.170 4.120 2.450 ;
        RECT  3.740 1.730 3.960 2.010 ;
        RECT  3.740 0.760 3.900 1.570 ;
        RECT  3.620 0.760 3.740 1.040 ;
        RECT  3.040 1.850 3.740 2.010 ;
        RECT  3.540 2.610 3.700 3.090 ;
        RECT  1.440 2.610 3.540 2.770 ;
        RECT  2.880 0.800 3.040 2.410 ;
        RECT  2.680 0.800 2.880 1.080 ;
        RECT  2.320 2.250 2.880 2.410 ;
        RECT  2.160 1.850 2.320 2.410 ;
        RECT  1.840 1.850 2.160 2.010 ;
        RECT  1.870 0.780 2.000 1.030 ;
        RECT  1.520 2.240 1.930 2.400 ;
        RECT  1.710 0.780 1.870 1.480 ;
        RECT  1.680 1.730 1.840 2.010 ;
        RECT  1.520 1.320 1.710 1.480 ;
        RECT  1.240 0.880 1.520 1.160 ;
        RECT  1.360 1.320 1.520 2.400 ;
        RECT  1.200 2.610 1.440 2.890 ;
        RECT  1.200 1.000 1.240 1.160 ;
        RECT  1.040 1.000 1.200 2.890 ;
        RECT  0.660 0.880 0.880 2.890 ;
    END
END MAS70

MACRO MAS71
    CLASS CORE ;
    FOREIGN MAS71 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.840 0.500 3.120 3.160 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 1.640 2.360 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.240 1.920 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.120 1.680 1.300 1.960 ;
        RECT  0.960 1.240 1.120 1.960 ;
        RECT  0.880 1.240 0.960 1.560 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.630 0.680 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 -0.280 3.200 0.280 ;
        RECT  2.220 -0.280 2.500 0.680 ;
        RECT  0.000 -0.280 2.220 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.580 3.320 3.200 3.880 ;
        RECT  2.300 2.440 2.580 3.880 ;
        RECT  1.540 3.260 2.300 3.880 ;
        RECT  1.260 2.440 1.540 3.880 ;
        RECT  0.540 3.260 1.260 3.880 ;
        RECT  0.260 2.230 0.540 3.880 ;
        RECT  0.000 3.320 0.260 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.520 0.920 2.680 2.280 ;
        RECT  0.880 0.920 2.520 1.080 ;
        RECT  2.060 2.120 2.520 2.280 ;
        RECT  1.780 2.120 2.060 2.400 ;
        RECT  1.020 2.120 1.780 2.280 ;
        RECT  0.740 2.120 1.020 2.400 ;
        RECT  0.600 0.800 0.880 1.080 ;
    END
END MAS71

MACRO MAS72
    CLASS CORE ;
    FOREIGN MAS72 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.950 0.520 2.110 3.160 ;
        RECT  1.650 0.520 1.950 0.780 ;
        RECT  1.500 2.840 1.950 3.160 ;
        END
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.270 2.840 2.720 3.160 ;
        END
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.850 1.060 2.130 ;
        RECT  0.480 1.850 0.760 2.360 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.240 3.120 2.360 ;
        RECT  2.840 1.240 2.880 1.730 ;
        RECT  2.650 1.450 2.840 1.730 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 -0.280 3.200 0.280 ;
        RECT  2.820 -0.280 3.110 0.740 ;
        RECT  0.930 -0.280 2.820 0.280 ;
        RECT  0.650 -0.280 0.930 1.290 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.110 3.320 3.200 3.880 ;
        RECT  2.880 2.770 3.110 3.880 ;
        RECT  0.940 3.320 2.880 3.880 ;
        RECT  0.660 2.960 0.940 3.880 ;
        RECT  0.000 3.320 0.660 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.490 1.010 2.550 1.290 ;
        RECT  2.270 1.010 2.490 2.550 ;
        RECT  1.630 0.960 1.790 2.530 ;
        RECT  1.370 0.960 1.630 1.120 ;
        RECT  1.340 2.370 1.630 2.530 ;
        RECT  1.250 1.530 1.470 1.960 ;
        RECT  1.210 0.460 1.370 1.120 ;
        RECT  1.060 2.370 1.340 2.650 ;
        RECT  0.370 1.530 1.250 1.690 ;
        RECT  1.090 0.460 1.210 0.740 ;
        RECT  0.320 1.010 0.370 1.690 ;
        RECT  0.160 1.010 0.320 2.550 ;
        RECT  0.090 1.010 0.160 1.290 ;
        RECT  0.090 2.270 0.160 2.550 ;
    END
END MAS72

MACRO MAS73
    CLASS CORE ;
    FOREIGN MAS73 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.930 0.800 1.240 1.080 ;
        RECT  0.690 0.920 0.930 1.080 ;
        RECT  0.690 2.040 0.920 2.410 ;
        RECT  0.530 0.920 0.690 2.410 ;
        RECT  0.480 2.040 0.530 2.410 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.530 0.370 1.810 ;
        RECT  0.080 1.530 0.320 2.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.850 1.240 1.160 1.660 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.370 -0.280 1.600 0.280 ;
        RECT  0.090 -0.280 0.370 1.310 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.440 3.320 1.600 3.880 ;
        RECT  1.180 2.030 1.440 3.880 ;
        RECT  0.380 3.260 1.180 3.880 ;
        RECT  0.140 2.920 0.380 3.880 ;
        RECT  0.000 3.320 0.140 3.880 ;
        END
    END VDD
END MAS73

MACRO MAS74
    CLASS CORE ;
    FOREIGN MAS74 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.440 1.120 2.430 ;
        RECT  0.870 0.440 0.880 1.230 ;
        RECT  0.680 2.120 0.880 2.430 ;
        RECT  0.680 0.840 0.870 1.230 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.680 1.640 0.720 1.960 ;
        RECT  0.400 1.390 0.680 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 -0.280 1.200 0.280 ;
        RECT  0.200 -0.280 0.480 1.220 ;
        RECT  0.000 -0.280 0.200 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 3.320 1.200 3.880 ;
        RECT  0.200 2.190 0.480 3.880 ;
        RECT  0.000 3.320 0.200 3.880 ;
        END
    END VDD
END MAS74

MACRO MAS75
    CLASS CORE ;
    FOREIGN MAS75 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.440 1.120 2.250 ;
        RECT  0.780 0.440 0.880 1.230 ;
        RECT  0.680 1.930 0.880 2.250 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.390 0.680 1.670 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 -0.280 1.200 0.280 ;
        RECT  0.160 -0.280 0.440 1.080 ;
        RECT  0.000 -0.280 0.160 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 3.320 1.200 3.880 ;
        RECT  0.160 2.520 0.440 3.880 ;
        RECT  0.000 3.320 0.160 3.880 ;
        END
    END VDD
END MAS75

MACRO MAS76
    CLASS CORE ;
    FOREIGN MAS76 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.840 2.320 2.280 ;
        RECT  0.890 0.920 2.080 1.080 ;
        RECT  1.810 2.120 2.080 2.280 ;
        RECT  1.530 2.120 1.810 2.550 ;
        END
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 0.840 0.510 1.480 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        RECT  0.480 1.640 0.880 1.960 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 1.920 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.520 1.960 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.090 -0.280 2.400 0.280 ;
        RECT  1.810 -0.280 2.090 0.350 ;
        RECT  0.370 -0.280 1.810 0.290 ;
        RECT  0.090 -0.280 0.370 0.370 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.850 3.320 2.400 3.880 ;
        RECT  0.570 2.440 0.850 3.880 ;
        RECT  0.000 3.320 0.570 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.170 2.440 2.290 2.690 ;
        RECT  2.010 2.440 2.170 3.100 ;
        RECT  1.330 2.940 2.010 3.100 ;
        RECT  1.170 2.120 1.330 3.100 ;
        RECT  1.050 2.120 1.170 2.550 ;
        RECT  0.370 2.120 1.050 2.280 ;
        RECT  0.090 2.120 0.370 2.580 ;
    END
END MAS76

MACRO MAS77
    CLASS CORE ;
    FOREIGN MAS77 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.110 0.440 1.120 1.560 ;
        RECT  0.950 0.440 1.110 3.100 ;
        RECT  0.880 0.440 0.950 1.560 ;
        RECT  0.790 2.400 0.950 3.100 ;
        RECT  0.800 0.840 0.880 1.160 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.450 1.580 0.720 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.550 -0.280 1.200 0.280 ;
        RECT  0.270 -0.280 0.550 1.250 ;
        RECT  0.000 -0.280 0.270 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.550 3.320 1.200 3.880 ;
        RECT  0.250 2.350 0.550 3.880 ;
        RECT  0.000 3.320 0.250 3.880 ;
        END
    END VDD
END MAS77

MACRO MAS78
    CLASS CORE ;
    FOREIGN MAS78 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.640 1.640 2.720 2.920 ;
        RECT  2.480 1.260 2.640 2.920 ;
        RECT  2.280 1.260 2.480 1.420 ;
        RECT  2.260 2.640 2.480 2.920 ;
        RECT  2.120 0.590 2.280 1.420 ;
        RECT  1.930 0.590 2.120 0.870 ;
        RECT  1.290 0.710 1.930 0.870 ;
        RECT  1.010 0.710 1.290 0.990 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.520 1.120 1.960 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.160 1.520 1.760 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.920 1.200 1.960 1.420 ;
        RECT  1.740 1.200 1.920 1.960 ;
        RECT  1.680 1.640 1.740 1.960 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.690 -0.280 2.800 0.280 ;
        RECT  2.440 -0.280 2.690 0.960 ;
        RECT  0.770 -0.280 2.440 0.280 ;
        RECT  0.490 -0.280 0.770 0.400 ;
        RECT  0.000 -0.280 0.490 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 3.320 2.800 3.880 ;
        RECT  0.760 2.840 1.040 3.880 ;
        RECT  0.000 3.320 0.760 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.080 1.580 2.300 2.280 ;
        RECT  1.880 2.120 2.080 2.280 ;
        RECT  1.720 2.120 1.880 2.680 ;
        RECT  0.680 2.490 1.720 2.680 ;
        RECT  0.520 0.920 0.680 2.680 ;
        RECT  0.370 0.920 0.520 1.080 ;
        RECT  0.210 2.520 0.520 2.680 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END MAS78

MACRO MAS79
    CLASS CORE ;
    FOREIGN MAS79 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.640 1.640 2.720 2.760 ;
        RECT  2.480 0.920 2.640 2.760 ;
        RECT  2.250 0.920 2.480 1.080 ;
        RECT  2.200 2.470 2.480 2.760 ;
        RECT  1.970 0.540 2.250 1.080 ;
        RECT  1.320 0.920 1.970 1.080 ;
        RECT  1.040 0.540 1.320 1.080 ;
        END
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.640 1.120 1.990 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.520 1.760 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.920 1.420 1.960 1.600 ;
        RECT  1.680 1.420 1.920 1.960 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.710 -0.280 2.800 0.280 ;
        RECT  2.430 -0.280 2.710 0.680 ;
        RECT  1.790 -0.280 2.430 0.280 ;
        RECT  1.510 -0.280 1.790 0.680 ;
        RECT  0.860 -0.280 1.510 0.280 ;
        RECT  0.580 -0.280 0.860 0.760 ;
        RECT  0.000 -0.280 0.580 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 3.320 2.800 3.880 ;
        RECT  0.800 2.470 1.040 3.880 ;
        RECT  0.000 3.320 0.800 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.080 1.760 2.320 2.310 ;
        RECT  0.640 2.150 2.080 2.310 ;
        RECT  0.480 0.920 0.640 2.690 ;
        RECT  0.370 0.920 0.480 1.080 ;
        RECT  0.210 2.530 0.480 2.690 ;
        RECT  0.090 0.800 0.370 1.080 ;
    END
END MAS79

MACRO MAS8
    CLASS CORE ;
    FOREIGN MAS8 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.440 1.920 2.610 ;
        RECT  1.680 0.440 1.760 1.560 ;
        RECT  1.390 2.450 1.760 2.610 ;
        RECT  1.640 0.840 1.680 1.160 ;
        RECT  1.080 2.450 1.390 2.680 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.160 1.920 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.520 0.720 1.960 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.020 -0.280 2.000 0.280 ;
        RECT  0.740 -0.280 1.020 0.400 ;
        RECT  0.000 -0.280 0.740 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.910 3.320 2.000 3.880 ;
        RECT  1.620 2.770 1.910 3.880 ;
        RECT  0.900 3.320 1.620 3.880 ;
        RECT  0.620 2.440 0.900 3.880 ;
        RECT  0.000 3.320 0.620 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.480 1.720 1.600 1.990 ;
        RECT  1.320 0.920 1.480 2.280 ;
        RECT  0.480 0.920 1.320 1.080 ;
        RECT  0.390 2.120 1.320 2.280 ;
        RECT  0.200 0.920 0.480 1.250 ;
        RECT  0.090 2.100 0.390 2.320 ;
    END
END MAS8

MACRO MAS80
    CLASS CORE ;
    FOREIGN MAS80 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.280 0.620 7.520 3.010 ;
        RECT  6.960 2.730 7.280 3.010 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.960 0.690 7.120 2.330 ;
        RECT  6.080 0.690 6.960 0.850 ;
        RECT  6.320 2.170 6.960 2.330 ;
        RECT  6.240 2.170 6.320 2.760 ;
        RECT  6.160 2.170 6.240 3.030 ;
        RECT  6.080 2.440 6.160 3.030 ;
        RECT  5.920 0.570 6.080 0.850 ;
        RECT  5.940 2.870 6.080 3.030 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 1.980 0.560 2.140 ;
        RECT  0.080 1.640 0.320 2.760 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.590 3.120 1.960 ;
        RECT  2.770 1.800 2.880 1.960 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.660 -0.280 7.600 0.280 ;
        RECT  6.380 -0.280 6.660 0.340 ;
        RECT  5.540 -0.280 6.380 0.280 ;
        RECT  5.260 -0.280 5.540 0.800 ;
        RECT  3.790 -0.280 5.260 0.280 ;
        RECT  3.510 -0.280 3.790 0.340 ;
        RECT  2.160 -0.280 3.510 0.280 ;
        RECT  2.000 -0.280 2.160 0.670 ;
        RECT  0.410 -0.280 2.000 0.280 ;
        RECT  0.130 -0.280 0.410 0.350 ;
        RECT  0.000 -0.280 0.130 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.640 3.320 7.600 3.880 ;
        RECT  6.480 2.490 6.640 3.880 ;
        RECT  5.360 3.320 6.480 3.880 ;
        RECT  5.080 2.860 5.360 3.880 ;
        RECT  3.660 3.320 5.080 3.880 ;
        RECT  3.380 3.260 3.660 3.880 ;
        RECT  2.550 3.320 3.380 3.880 ;
        RECT  1.870 3.260 2.550 3.880 ;
        RECT  0.410 3.320 1.870 3.880 ;
        RECT  0.130 3.260 0.410 3.880 ;
        RECT  0.000 3.320 0.130 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  6.570 1.090 6.800 2.010 ;
        RECT  5.820 1.090 6.570 1.250 ;
        RECT  5.820 1.850 6.570 2.010 ;
        RECT  5.670 1.410 6.240 1.690 ;
        RECT  5.660 1.850 5.820 2.630 ;
        RECT  4.980 1.410 5.670 1.570 ;
        RECT  5.420 1.850 5.660 2.010 ;
        RECT  5.140 1.740 5.420 2.010 ;
        RECT  4.820 0.840 4.980 2.420 ;
        RECT  4.270 0.840 4.820 1.000 ;
        RECT  4.440 2.260 4.820 2.420 ;
        RECT  4.500 1.160 4.660 2.100 ;
        RECT  3.760 1.160 4.500 1.320 ;
        RECT  4.120 1.940 4.500 2.100 ;
        RECT  4.280 2.260 4.440 3.010 ;
        RECT  3.440 1.540 4.310 1.700 ;
        RECT  3.960 1.940 4.120 3.070 ;
        RECT  1.530 2.910 3.960 3.070 ;
        RECT  3.640 1.880 3.800 2.750 ;
        RECT  3.600 0.640 3.760 1.320 ;
        RECT  2.490 2.590 3.640 2.750 ;
        RECT  2.870 0.640 3.600 0.800 ;
        RECT  3.280 1.150 3.440 2.430 ;
        RECT  3.160 1.150 3.280 1.310 ;
        RECT  2.940 2.270 3.280 2.430 ;
        RECT  3.000 0.960 3.160 1.310 ;
        RECT  1.840 0.960 3.000 1.120 ;
        RECT  2.710 0.510 2.870 0.800 ;
        RECT  2.590 0.510 2.710 0.670 ;
        RECT  2.490 1.280 2.610 2.260 ;
        RECT  2.450 1.280 2.490 2.750 ;
        RECT  2.330 1.280 2.450 1.440 ;
        RECT  2.330 2.100 2.450 2.750 ;
        RECT  1.850 2.100 2.330 2.260 ;
        RECT  2.130 1.600 2.290 1.940 ;
        RECT  1.520 1.600 2.130 1.760 ;
        RECT  1.690 1.920 1.850 2.260 ;
        RECT  1.680 0.450 1.840 1.120 ;
        RECT  1.220 0.450 1.680 0.610 ;
        RECT  1.370 1.980 1.530 3.070 ;
        RECT  1.360 0.850 1.520 1.760 ;
        RECT  1.200 1.980 1.370 2.140 ;
        RECT  0.650 0.850 1.360 1.010 ;
        RECT  1.050 2.300 1.210 2.580 ;
        RECT  1.040 1.200 1.200 2.140 ;
        RECT  0.880 2.300 1.050 2.460 ;
        RECT  0.820 1.200 1.040 1.480 ;
        RECT  0.720 1.660 0.880 2.460 ;
        RECT  0.650 1.660 0.720 1.820 ;
        RECT  0.490 0.850 0.650 1.820 ;
    END
END MAS80

MACRO MAS81
    CLASS CORE ;
    FOREIGN MAS81 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.840 1.030 7.120 2.360 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.520 0.560 6.680 2.200 ;
        RECT  5.940 0.560 6.520 0.720 ;
        RECT  6.360 2.040 6.520 2.200 ;
        RECT  6.240 2.040 6.360 2.360 ;
        RECT  6.080 2.040 6.240 3.070 ;
        RECT  5.700 2.790 6.080 3.070 ;
        RECT  5.660 0.440 5.940 0.720 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.430 2.440 0.720 2.760 ;
        RECT  0.270 1.960 0.430 2.760 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  2.840 1.590 3.120 1.960 ;
        RECT  2.770 1.680 2.840 1.960 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 -0.280 7.200 0.280 ;
        RECT  6.220 -0.280 6.500 0.400 ;
        RECT  5.480 -0.280 6.220 0.280 ;
        RECT  5.200 -0.280 5.480 0.400 ;
        RECT  3.480 -0.280 5.200 0.340 ;
        RECT  2.210 -0.280 3.480 0.280 ;
        RECT  1.930 -0.280 2.210 0.670 ;
        RECT  0.400 -0.280 1.930 0.340 ;
        RECT  0.120 -0.280 0.400 0.400 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  6.680 3.320 7.200 3.880 ;
        RECT  6.400 2.640 6.680 3.880 ;
        RECT  5.360 3.320 6.400 3.880 ;
        RECT  5.080 2.710 5.360 3.880 ;
        RECT  3.360 3.260 5.080 3.880 ;
        RECT  2.490 3.320 3.360 3.880 ;
        RECT  1.810 3.260 2.490 3.880 ;
        RECT  0.400 3.320 1.810 3.880 ;
        RECT  0.120 3.200 0.400 3.880 ;
        RECT  0.000 3.320 0.120 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  6.240 1.580 6.360 1.880 ;
        RECT  6.080 0.900 6.240 1.880 ;
        RECT  5.660 0.900 6.080 1.120 ;
        RECT  5.800 1.720 6.080 1.880 ;
        RECT  5.640 1.280 5.920 1.560 ;
        RECT  5.800 2.270 5.920 2.550 ;
        RECT  5.640 1.720 5.800 2.550 ;
        RECT  5.040 1.280 5.640 1.440 ;
        RECT  5.480 1.720 5.640 1.880 ;
        RECT  5.200 1.600 5.480 1.880 ;
        RECT  4.880 0.590 5.040 2.390 ;
        RECT  4.240 0.590 4.880 0.870 ;
        RECT  4.580 2.230 4.880 2.390 ;
        RECT  4.440 1.030 4.720 1.950 ;
        RECT  4.360 2.230 4.580 2.510 ;
        RECT  3.760 1.030 4.440 1.190 ;
        RECT  4.320 1.790 4.440 1.950 ;
        RECT  4.200 1.790 4.320 2.070 ;
        RECT  4.000 1.350 4.280 1.630 ;
        RECT  4.040 1.790 4.200 3.100 ;
        RECT  1.530 2.880 4.040 3.100 ;
        RECT  3.440 1.350 4.000 1.510 ;
        RECT  3.600 1.790 3.880 2.720 ;
        RECT  3.600 0.500 3.760 1.190 ;
        RECT  2.840 0.500 3.600 0.780 ;
        RECT  2.530 2.560 3.600 2.720 ;
        RECT  3.280 1.060 3.440 2.400 ;
        RECT  3.190 1.060 3.280 1.220 ;
        RECT  2.910 2.120 3.280 2.400 ;
        RECT  2.910 0.940 3.190 1.220 ;
        RECT  1.770 0.940 2.910 1.100 ;
        RECT  2.680 0.450 2.840 0.780 ;
        RECT  2.560 0.450 2.680 0.670 ;
        RECT  2.530 1.260 2.610 2.240 ;
        RECT  2.450 1.260 2.530 2.720 ;
        RECT  2.330 1.260 2.450 1.480 ;
        RECT  2.250 2.080 2.450 2.720 ;
        RECT  2.170 1.640 2.290 1.920 ;
        RECT  1.850 2.080 2.250 2.240 ;
        RECT  2.010 1.260 2.170 1.920 ;
        RECT  1.450 1.260 2.010 1.420 ;
        RECT  1.570 1.960 1.850 2.240 ;
        RECT  1.610 0.500 1.770 1.100 ;
        RECT  1.120 0.500 1.610 0.720 ;
        RECT  1.390 2.400 1.530 3.100 ;
        RECT  1.290 0.880 1.450 1.420 ;
        RECT  1.370 1.580 1.390 3.100 ;
        RECT  1.230 1.580 1.370 2.560 ;
        RECT  0.450 0.880 1.290 1.100 ;
        RECT  1.130 1.580 1.230 1.740 ;
        RECT  1.050 2.880 1.210 3.160 ;
        RECT  0.970 1.260 1.130 1.740 ;
        RECT  0.890 1.900 1.050 3.160 ;
        RECT  0.640 1.260 0.970 1.480 ;
        RECT  0.810 1.900 0.890 2.060 ;
        RECT  0.650 1.640 0.810 2.060 ;
        RECT  0.450 1.640 0.650 1.800 ;
        RECT  0.290 0.880 0.450 1.800 ;
    END
END MAS81

MACRO MAS82
    CLASS CORE ;
    FOREIGN MAS82 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.210 0.440 2.320 1.560 ;
        RECT  2.080 0.440 2.210 2.350 ;
        RECT  1.930 0.520 2.080 2.350 ;
        RECT  1.130 0.520 1.930 0.760 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.800 1.360 1.120 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.600 1.680 ;
        END
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.940 -0.280 2.400 0.280 ;
        RECT  0.670 -0.280 0.940 0.750 ;
        RECT  0.000 -0.280 0.670 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.050 3.320 2.400 3.880 ;
        RECT  0.770 2.840 1.050 3.880 ;
        RECT  0.000 3.320 0.770 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.370 2.660 2.010 2.940 ;
        RECT  1.210 2.520 1.370 2.940 ;
        RECT  0.640 2.520 1.210 2.680 ;
        RECT  0.480 0.920 0.640 2.680 ;
        RECT  0.090 0.920 0.480 1.080 ;
        RECT  0.370 2.520 0.480 2.680 ;
        RECT  0.090 2.520 0.370 2.800 ;
    END
END MAS82

MACRO MAS83
    CLASS CORE ;
    FOREIGN MAS83 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 1.240 1.920 2.360 ;
        RECT  1.680 0.920 1.760 2.360 ;
        RECT  1.600 0.920 1.680 2.300 ;
        RECT  1.300 0.920 1.600 1.080 ;
        RECT  1.190 2.120 1.600 2.300 ;
        RECT  1.020 0.440 1.300 1.080 ;
        RECT  0.910 2.120 1.190 2.870 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.440 1.640 ;
        RECT  0.720 1.240 1.280 1.400 ;
        RECT  0.540 1.240 0.720 1.560 ;
        RECT  0.310 1.240 0.540 1.870 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.640 1.120 1.960 ;
        RECT  0.800 1.740 0.880 1.960 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.820 -0.280 2.000 0.280 ;
        RECT  1.540 -0.280 1.820 0.760 ;
        RECT  0.830 -0.280 1.540 0.280 ;
        RECT  0.530 -0.280 0.830 1.080 ;
        RECT  0.000 -0.280 0.530 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.880 3.320 2.000 3.880 ;
        RECT  1.640 3.220 1.880 3.880 ;
        RECT  0.410 3.320 1.640 3.880 ;
        RECT  0.110 2.150 0.410 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
END MAS83

MACRO MAS84
    CLASS CORE ;
    FOREIGN MAS84 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.940 0.800 1.120 2.160 ;
        RECT  0.880 0.800 0.940 3.020 ;
        RECT  0.660 0.800 0.880 1.080 ;
        RECT  0.660 1.910 0.880 3.020 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.240 0.720 1.630 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.450 -0.280 1.600 0.280 ;
        RECT  1.280 -0.280 1.450 1.060 ;
        RECT  0.420 -0.280 1.280 0.340 ;
        RECT  0.140 -0.280 0.420 1.080 ;
        RECT  0.000 -0.280 0.140 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.460 3.320 1.600 3.880 ;
        RECT  1.180 2.400 1.460 3.880 ;
        RECT  0.460 3.320 1.180 3.880 ;
        RECT  0.180 1.910 0.460 3.880 ;
        RECT  0.000 3.320 0.180 3.880 ;
        END
    END VDD
END MAS84

MACRO MAS85
    CLASS CORE ;
    FOREIGN MAS85 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.700 1.560 4.720 2.760 ;
        RECT  4.420 0.600 4.700 2.760 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.670 4.260 2.600 ;
        RECT  3.700 0.670 4.100 0.830 ;
        RECT  3.560 2.440 4.100 2.600 ;
        RECT  3.420 0.550 3.700 0.830 ;
        RECT  3.270 2.440 3.560 2.950 ;
        END
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.500 0.430 1.780 ;
        RECT  0.320 1.500 0.360 1.960 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.380 1.220 1.960 1.600 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.290 -0.280 4.800 0.280 ;
        RECT  4.010 -0.280 4.290 0.360 ;
        RECT  3.160 -0.280 4.010 0.280 ;
        RECT  2.920 -0.280 3.160 0.820 ;
        RECT  1.420 -0.280 2.920 0.280 ;
        RECT  1.120 -0.280 1.420 0.590 ;
        RECT  0.370 -0.280 1.120 0.280 ;
        RECT  0.090 -0.280 0.370 0.640 ;
        RECT  0.000 -0.280 0.090 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  4.170 3.320 4.800 3.880 ;
        RECT  3.840 2.910 4.170 3.880 ;
        RECT  3.080 3.320 3.840 3.880 ;
        RECT  2.780 2.800 3.080 3.880 ;
        RECT  1.540 3.320 2.780 3.880 ;
        RECT  1.260 2.930 1.540 3.880 ;
        RECT  0.370 3.320 1.260 3.880 ;
        RECT  0.090 3.240 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  3.700 1.410 3.940 1.690 ;
        RECT  3.580 1.010 3.700 1.690 ;
        RECT  3.420 1.010 3.580 2.270 ;
        RECT  2.820 1.990 3.420 2.270 ;
        RECT  3.040 1.380 3.260 1.660 ;
        RECT  2.760 1.380 3.040 1.540 ;
        RECT  2.660 1.720 2.820 2.270 ;
        RECT  2.600 0.580 2.760 1.540 ;
        RECT  2.540 1.720 2.660 1.940 ;
        RECT  2.260 0.580 2.600 0.740 ;
        RECT  2.280 1.340 2.600 1.540 ;
        RECT  2.220 0.900 2.440 1.180 ;
        RECT  2.120 1.340 2.280 2.170 ;
        RECT  1.980 0.460 2.260 0.740 ;
        RECT  1.220 0.900 2.220 1.060 ;
        RECT  1.900 1.890 2.120 2.170 ;
        RECT  1.860 2.660 1.980 2.940 ;
        RECT  1.700 2.540 1.860 2.940 ;
        RECT  1.220 2.540 1.700 2.750 ;
        RECT  1.060 0.750 1.220 2.750 ;
        RECT  0.820 2.920 1.100 3.160 ;
        RECT  0.830 0.750 1.060 0.910 ;
        RECT  0.620 2.480 1.060 2.750 ;
        RECT  0.620 1.070 0.900 2.290 ;
        RECT  0.550 0.550 0.830 0.910 ;
        RECT  0.420 2.920 0.820 3.080 ;
        RECT  0.530 1.070 0.620 1.290 ;
        RECT  0.510 2.030 0.620 2.290 ;
        RECT  0.420 2.130 0.510 2.290 ;
        RECT  0.260 2.130 0.420 3.080 ;
    END
END MAS85

MACRO MAS86
    CLASS CORE ;
    FOREIGN MAS86 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.220 1.520 1.700 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.080 0.500 8.320 2.890 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.280 1.090 7.520 2.270 ;
        RECT  7.040 1.090 7.280 1.310 ;
        RECT  7.040 1.910 7.280 2.270 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.960 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  2.040 1.220 2.320 1.560 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.800 -0.280 8.400 0.280 ;
        RECT  7.520 -0.280 7.800 0.610 ;
        RECT  6.400 -0.280 7.520 0.280 ;
        RECT  5.920 -0.280 6.400 0.400 ;
        RECT  4.300 -0.280 5.920 0.340 ;
        RECT  4.020 -0.280 4.300 0.990 ;
        RECT  2.520 -0.280 4.020 0.340 ;
        RECT  2.240 -0.280 2.520 0.400 ;
        RECT  1.620 -0.280 2.240 0.280 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  0.730 -0.280 1.340 0.340 ;
        RECT  0.000 -0.280 0.730 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  7.800 3.320 8.400 3.880 ;
        RECT  7.520 2.990 7.800 3.880 ;
        RECT  6.370 3.320 7.520 3.880 ;
        RECT  6.090 2.850 6.370 3.880 ;
        RECT  4.000 3.260 6.090 3.880 ;
        RECT  3.720 2.400 4.000 3.880 ;
        RECT  2.520 3.260 3.720 3.880 ;
        RECT  2.240 3.210 2.520 3.880 ;
        RECT  1.400 3.320 2.240 3.880 ;
        RECT  1.120 3.210 1.400 3.880 ;
        RECT  0.470 3.260 1.120 3.880 ;
        RECT  0.000 3.320 0.470 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  7.760 0.770 7.920 2.810 ;
        RECT  6.960 0.770 7.760 0.930 ;
        RECT  6.920 2.650 7.760 2.810 ;
        RECT  6.640 1.560 7.120 1.720 ;
        RECT  6.680 0.450 6.960 0.930 ;
        RECT  6.760 2.650 6.920 3.150 ;
        RECT  6.580 2.910 6.760 3.150 ;
        RECT  6.600 1.090 6.640 1.720 ;
        RECT  6.440 1.090 6.600 2.600 ;
        RECT  6.360 1.090 6.440 1.720 ;
        RECT  6.300 2.340 6.440 2.600 ;
        RECT  5.680 1.560 6.360 1.720 ;
        RECT  5.320 1.900 6.280 2.180 ;
        RECT  5.220 2.710 5.500 2.990 ;
        RECT  5.260 0.920 5.320 2.180 ;
        RECT  5.040 0.920 5.260 2.500 ;
        RECT  4.400 2.710 5.220 2.870 ;
        RECT  4.980 2.220 5.040 2.500 ;
        RECT  4.720 0.730 4.860 1.010 ;
        RECT  4.560 0.730 4.720 2.540 ;
        RECT  4.180 1.150 4.560 1.310 ;
        RECT  4.240 1.590 4.400 2.870 ;
        RECT  3.680 1.590 4.240 1.750 ;
        RECT  3.900 1.150 4.180 1.430 ;
        RECT  3.420 1.910 4.080 2.190 ;
        RECT  3.520 0.500 3.680 1.750 ;
        RECT  3.040 0.500 3.520 0.780 ;
        RECT  3.360 1.910 3.420 2.680 ;
        RECT  3.200 1.030 3.360 2.680 ;
        RECT  2.960 2.440 3.200 2.680 ;
        RECT  2.940 0.500 3.040 2.280 ;
        RECT  2.800 2.440 2.960 3.050 ;
        RECT  2.880 0.570 2.940 2.280 ;
        RECT  2.800 0.570 2.880 0.850 ;
        RECT  2.800 1.910 2.880 2.280 ;
        RECT  0.680 2.120 2.800 2.280 ;
        RECT  0.370 2.890 2.800 3.050 ;
        RECT  2.640 1.220 2.720 1.500 ;
        RECT  2.480 0.900 2.640 1.940 ;
        RECT  2.080 0.900 2.480 1.060 ;
        RECT  1.680 1.720 2.480 1.940 ;
        RECT  1.800 0.780 2.080 1.060 ;
        RECT  0.600 2.460 1.920 2.730 ;
        RECT  0.800 0.900 1.800 1.060 ;
        RECT  0.640 0.500 0.800 1.060 ;
        RECT  0.400 1.980 0.680 2.280 ;
        RECT  0.440 0.500 0.640 0.780 ;
        RECT  0.240 0.940 0.480 1.220 ;
        RECT  0.240 2.440 0.370 3.050 ;
        RECT  0.210 0.940 0.240 3.050 ;
        RECT  0.080 0.940 0.210 2.720 ;
    END
END MAS86

MACRO MAS87
    CLASS CORE ;
    FOREIGN MAS87 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.360 1.040 2.730 1.760 ;
        RECT  2.280 1.040 2.360 3.160 ;
        RECT  2.110 0.600 2.280 3.160 ;
        RECT  2.040 0.600 2.110 1.280 ;
        RECT  2.080 2.020 2.110 3.160 ;
        RECT  1.920 0.600 2.040 0.760 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.560 1.750 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.520 1.120 1.960 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.420 1.240 0.720 1.670 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.710 -0.280 3.200 0.280 ;
        RECT  2.440 -0.280 2.710 0.820 ;
        RECT  1.720 -0.280 2.440 0.280 ;
        RECT  1.440 -0.280 1.720 0.650 ;
        RECT  0.000 -0.280 1.440 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.920 3.320 3.200 3.880 ;
        RECT  2.640 2.020 2.920 3.880 ;
        RECT  1.880 3.320 2.640 3.880 ;
        RECT  1.600 2.440 1.880 3.880 ;
        RECT  0.920 3.320 1.600 3.880 ;
        RECT  0.640 2.440 0.920 3.880 ;
        RECT  0.000 3.320 0.640 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.880 1.490 1.940 1.770 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  0.520 0.920 1.720 1.080 ;
        RECT  1.400 2.120 1.720 2.280 ;
        RECT  1.120 2.120 1.400 2.950 ;
        RECT  0.440 2.120 1.120 2.280 ;
        RECT  0.240 0.740 0.520 1.080 ;
        RECT  0.160 2.120 0.440 2.950 ;
    END
END MAS87

MACRO MAS88
    CLASS CORE ;
    FOREIGN MAS88 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.060 1.640 3.220 1.960 ;
        RECT  2.880 1.600 3.060 1.960 ;
        END
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.650 0.840 9.920 2.650 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.430 1.240 2.720 1.560 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.240 0.760 1.640 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  3.740 -0.280 10.000 0.280 ;
        RECT  2.120 -0.280 3.740 0.340 ;
        RECT  0.930 -0.280 2.120 0.280 ;
        RECT  0.650 -0.280 0.930 0.400 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  9.390 3.320 10.000 3.880 ;
        RECT  8.450 2.770 9.390 3.880 ;
        RECT  6.410 3.320 8.450 3.880 ;
        RECT  5.100 3.260 6.410 3.880 ;
        RECT  3.860 3.320 5.100 3.880 ;
        RECT  3.580 3.200 3.860 3.880 ;
        RECT  2.400 3.320 3.580 3.880 ;
        RECT  2.120 3.200 2.400 3.880 ;
        RECT  0.810 3.260 2.120 3.880 ;
        RECT  0.530 2.800 0.810 3.880 ;
        RECT  0.000 3.320 0.530 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  9.310 1.300 9.430 1.580 ;
        RECT  9.150 0.440 9.310 2.510 ;
        RECT  7.390 0.440 9.150 0.660 ;
        RECT  7.430 2.350 9.150 2.510 ;
        RECT  8.830 1.030 8.950 1.310 ;
        RECT  8.830 1.910 8.950 2.190 ;
        RECT  8.670 1.030 8.830 2.190 ;
        RECT  8.290 1.350 8.670 1.630 ;
        RECT  8.230 0.820 8.510 1.100 ;
        RECT  8.130 0.940 8.230 1.100 ;
        RECT  8.010 0.940 8.130 1.820 ;
        RECT  7.970 0.940 8.010 2.190 ;
        RECT  7.850 1.540 7.970 2.190 ;
        RECT  7.310 2.030 7.850 2.190 ;
        RECT  6.570 2.940 7.760 3.160 ;
        RECT  7.470 0.820 7.690 1.870 ;
        RECT  7.230 0.820 7.470 0.980 ;
        RECT  7.150 2.350 7.430 2.630 ;
        RECT  7.150 1.140 7.310 2.190 ;
        RECT  7.070 0.440 7.230 0.980 ;
        RECT  6.910 1.140 7.150 1.300 ;
        RECT  4.060 0.440 7.070 0.600 ;
        RECT  6.830 1.460 6.990 2.500 ;
        RECT  6.750 0.760 6.910 1.300 ;
        RECT  6.590 1.460 6.830 1.620 ;
        RECT  6.240 2.220 6.830 2.500 ;
        RECT  4.380 0.760 6.750 0.920 ;
        RECT  6.450 1.780 6.670 2.060 ;
        RECT  6.310 1.080 6.590 1.620 ;
        RECT  4.940 2.940 6.570 3.100 ;
        RECT  5.800 1.780 6.450 1.940 ;
        RECT  6.080 2.100 6.240 2.500 ;
        RECT  5.960 2.100 6.080 2.380 ;
        RECT  5.640 1.140 5.800 2.780 ;
        RECT  4.940 1.140 5.640 1.300 ;
        RECT  5.320 2.500 5.640 2.780 ;
        RECT  4.940 2.060 5.480 2.340 ;
        RECT  4.660 1.080 4.940 1.300 ;
        RECT  4.780 1.520 4.940 3.100 ;
        RECT  4.300 1.520 4.780 1.680 ;
        RECT  4.180 2.940 4.780 3.100 ;
        RECT  3.860 1.140 4.660 1.300 ;
        RECT  4.400 2.500 4.620 2.780 ;
        RECT  3.860 1.910 4.420 2.190 ;
        RECT  3.100 2.500 4.400 2.660 ;
        RECT  4.220 0.760 4.380 0.980 ;
        RECT  4.020 1.460 4.300 1.680 ;
        RECT  3.540 0.820 4.220 0.980 ;
        RECT  4.020 2.880 4.180 3.100 ;
        RECT  3.900 0.440 4.060 0.660 ;
        RECT  3.420 2.880 4.020 3.040 ;
        RECT  1.840 0.500 3.900 0.660 ;
        RECT  3.700 1.140 3.860 2.190 ;
        RECT  3.380 0.820 3.540 2.280 ;
        RECT  3.260 2.880 3.420 3.130 ;
        RECT  3.020 0.820 3.380 1.040 ;
        RECT  3.020 2.120 3.380 2.280 ;
        RECT  2.720 2.970 3.260 3.130 ;
        RECT  2.880 2.500 3.100 2.810 ;
        RECT  2.510 2.500 2.880 2.660 ;
        RECT  2.270 0.820 2.840 1.040 ;
        RECT  2.560 2.820 2.720 3.130 ;
        RECT  1.730 2.820 2.560 2.980 ;
        RECT  2.350 1.740 2.510 2.660 ;
        RECT  2.270 1.740 2.350 1.900 ;
        RECT  2.110 0.820 2.270 1.900 ;
        RECT  1.910 2.060 2.190 2.340 ;
        RECT  1.840 2.060 1.910 2.220 ;
        RECT  1.680 0.500 1.840 2.220 ;
        RECT  1.570 2.380 1.730 2.980 ;
        RECT  1.560 0.500 1.680 0.960 ;
        RECT  1.250 1.760 1.680 2.040 ;
        RECT  1.450 2.380 1.570 2.660 ;
        RECT  1.090 2.380 1.450 2.540 ;
        RECT  1.120 0.440 1.400 0.720 ;
        RECT  1.090 1.030 1.370 1.310 ;
        RECT  0.310 0.560 1.120 0.720 ;
        RECT  0.930 1.030 1.090 2.540 ;
        RECT  0.150 0.560 0.310 2.320 ;
    END
END MAS88

MACRO MAS89
    CLASS CORE ;
    FOREIGN MAS89 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 1.210 2.320 1.570 ;
        RECT  1.890 0.970 2.180 2.490 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 0.840 1.120 1.380 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.320 2.820 0.720 3.160 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.800 -0.280 3.200 0.280 ;
        RECT  0.930 -0.280 2.800 0.340 ;
        RECT  0.650 -0.280 0.930 0.680 ;
        RECT  0.000 -0.280 0.650 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.730 3.320 3.200 3.880 ;
        RECT  2.450 3.200 2.730 3.880 ;
        RECT  1.050 3.260 2.450 3.880 ;
        RECT  0.880 2.330 1.050 3.880 ;
        RECT  0.770 2.330 0.880 2.620 ;
        RECT  0.000 3.320 0.880 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  2.960 0.630 3.120 1.710 ;
        RECT  1.730 0.630 2.960 0.790 ;
        RECT  2.840 1.430 2.960 1.710 ;
        RECT  2.680 0.950 2.800 1.230 ;
        RECT  2.680 2.210 2.800 3.000 ;
        RECT  2.520 0.950 2.680 3.000 ;
        RECT  1.570 0.630 1.730 2.370 ;
        RECT  1.310 0.770 1.570 1.050 ;
        RECT  1.530 2.210 1.570 2.370 ;
        RECT  1.250 2.210 1.530 2.490 ;
        RECT  1.130 1.540 1.410 1.820 ;
        RECT  0.370 1.660 1.130 1.820 ;
        RECT  0.210 0.850 0.370 2.490 ;
        RECT  0.090 0.850 0.210 1.130 ;
        RECT  0.090 2.210 0.210 2.490 ;
    END
END MAS89

MACRO MAS9
    CLASS CORE ;
    FOREIGN MAS9 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.110 0.530 6.320 3.160 ;
        RECT  6.090 0.530 6.110 0.840 ;
        RECT  6.080 1.910 6.110 3.160 ;
        END
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 0.440 4.360 0.760 ;
        END
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 2.840 1.140 3.160 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.840 0.320 1.960 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.240 1.720 1.640 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 1.520 3.560 1.960 ;
        RECT  3.220 1.520 3.280 1.800 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  5.790 -0.280 6.400 0.280 ;
        RECT  5.510 -0.280 5.790 0.510 ;
        RECT  3.600 -0.280 5.510 0.280 ;
        RECT  3.280 -0.280 3.600 0.870 ;
        RECT  1.560 -0.280 3.280 0.340 ;
        RECT  1.280 -0.280 1.560 1.030 ;
        RECT  0.380 -0.280 1.280 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        RECT  0.000 -0.280 0.100 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  5.900 3.320 6.400 3.880 ;
        RECT  5.620 3.000 5.900 3.880 ;
        RECT  3.640 3.320 5.620 3.880 ;
        RECT  3.360 3.260 3.640 3.880 ;
        RECT  1.520 3.320 3.360 3.880 ;
        RECT  1.300 2.780 1.520 3.880 ;
        RECT  0.380 3.320 1.300 3.880 ;
        RECT  0.100 3.200 0.380 3.880 ;
        RECT  0.000 3.320 0.100 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  5.870 1.370 5.950 1.650 ;
        RECT  5.710 0.670 5.870 1.650 ;
        RECT  5.080 0.670 5.710 0.830 ;
        RECT  5.520 1.030 5.550 1.420 ;
        RECT  5.400 1.030 5.520 2.530 ;
        RECT  5.360 1.030 5.400 3.100 ;
        RECT  5.220 2.250 5.360 3.100 ;
        RECT  1.840 2.940 5.220 3.100 ;
        RECT  4.960 0.670 5.080 1.220 ;
        RECT  4.800 0.670 4.960 2.440 ;
        RECT  4.680 2.160 4.800 2.440 ;
        RECT  4.480 0.960 4.640 2.000 ;
        RECT  4.320 0.960 4.480 1.240 ;
        RECT  4.320 1.840 4.480 2.780 ;
        RECT  4.140 1.400 4.320 1.680 ;
        RECT  2.740 2.560 4.320 2.780 ;
        RECT  3.860 0.920 4.140 2.360 ;
        RECT  3.060 2.080 3.120 2.360 ;
        RECT  2.900 0.620 3.060 2.360 ;
        RECT  2.780 0.620 2.900 0.900 ;
        RECT  2.580 1.060 2.740 2.780 ;
        RECT  2.520 1.060 2.580 1.220 ;
        RECT  2.240 2.500 2.580 2.780 ;
        RECT  2.240 0.820 2.520 1.220 ;
        RECT  2.260 1.380 2.420 2.300 ;
        RECT  2.040 1.380 2.260 1.540 ;
        RECT  1.760 2.140 2.260 2.300 ;
        RECT  1.880 1.700 2.100 1.980 ;
        RECT  1.880 0.800 2.040 1.540 ;
        RECT  1.760 0.800 1.880 1.080 ;
        RECT  1.120 1.820 1.880 1.980 ;
        RECT  1.680 2.460 1.840 3.100 ;
        RECT  0.800 2.460 1.680 2.620 ;
        RECT  0.960 0.490 1.120 2.220 ;
        RECT  0.720 0.490 0.960 0.770 ;
        RECT  0.840 1.940 0.960 2.220 ;
        RECT  0.680 1.030 0.800 1.310 ;
        RECT  0.680 2.460 0.800 2.680 ;
        RECT  0.520 1.030 0.680 2.680 ;
    END
END MAS9

MACRO MAS90
    CLASS CORE ;
    FOREIGN MAS90 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.580 0.840 4.720 2.070 ;
        RECT  4.360 0.440 4.580 3.160 ;
        RECT  4.300 0.440 4.360 1.340 ;
        RECT  4.300 1.880 4.360 3.160 ;
        END
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 1.640 2.400 2.360 ;
        RECT  2.080 2.040 2.240 2.360 ;
        END
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.880 1.640 3.350 1.960 ;
        END
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.240 0.320 2.360 ;
        END
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.150 0.890 1.560 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.920 1.640 2.070 1.880 ;
        RECT  1.680 1.640 1.920 2.070 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 1.800 1.520 2.360 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  5.060 -0.280 5.200 0.280 ;
        RECT  4.780 -0.280 5.060 0.670 ;
        RECT  4.060 -0.280 4.780 0.280 ;
        RECT  0.120 -0.280 4.060 0.340 ;
        RECT  0.000 -0.280 0.120 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  5.060 3.320 5.200 3.880 ;
        RECT  4.780 2.230 5.060 3.880 ;
        RECT  4.100 3.320 4.780 3.880 ;
        RECT  3.820 2.440 4.100 3.880 ;
        RECT  2.250 3.260 3.820 3.880 ;
        RECT  1.970 3.200 2.250 3.880 ;
        RECT  0.610 3.260 1.970 3.880 ;
        RECT  0.330 2.610 0.610 3.880 ;
        RECT  0.000 3.320 0.330 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  4.080 1.470 4.180 1.750 ;
        RECT  3.920 1.000 4.080 2.280 ;
        RECT  3.620 1.000 3.920 1.160 ;
        RECT  3.620 2.120 3.920 2.280 ;
        RECT  3.540 1.320 3.760 1.660 ;
        RECT  3.340 0.880 3.620 1.160 ;
        RECT  3.340 2.120 3.620 3.100 ;
        RECT  2.760 1.320 3.540 1.480 ;
        RECT  2.810 2.520 3.090 2.800 ;
        RECT  2.720 2.520 2.810 2.680 ;
        RECT  2.720 1.200 2.760 1.480 ;
        RECT  2.560 1.200 2.720 2.680 ;
        RECT  2.480 1.200 2.560 1.480 ;
        RECT  1.410 2.520 2.560 2.680 ;
        RECT  2.000 1.170 2.280 1.450 ;
        RECT  1.360 1.290 2.000 1.450 ;
        RECT  1.480 0.700 1.760 0.980 ;
        RECT  0.830 0.820 1.480 0.980 ;
        RECT  1.130 2.520 1.410 2.800 ;
        RECT  1.070 1.290 1.360 1.570 ;
        RECT  0.610 0.700 0.830 0.980 ;
    END
END MAS90

MACRO MAS91
    CLASS CORE ;
    FOREIGN MAS91 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.430 1.360 6.690 1.640 ;
        RECT  6.050 1.360 6.430 1.520 ;
        RECT  5.890 0.470 6.050 1.520 ;
        RECT  4.810 0.470 5.890 0.630 ;
        RECT  4.650 0.470 4.810 1.010 ;
        RECT  4.490 0.850 4.650 1.010 ;
        RECT  4.210 0.850 4.490 1.510 ;
        RECT  4.170 0.850 4.210 1.010 ;
        RECT  4.010 0.440 4.170 1.010 ;
        RECT  1.900 0.440 4.010 0.600 ;
        RECT  1.740 0.440 1.900 0.700 ;
        RECT  1.120 0.540 1.740 0.700 ;
        RECT  1.200 1.360 1.440 1.640 ;
        RECT  1.120 1.360 1.200 1.560 ;
        RECT  0.960 0.540 1.120 1.560 ;
        RECT  0.880 0.840 0.960 1.560 ;
        END
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.270 1.640 8.320 2.390 ;
        RECT  8.150 1.150 8.270 2.390 ;
        RECT  8.110 1.030 8.150 2.390 ;
        RECT  7.830 1.030 8.110 1.310 ;
        RECT  8.080 1.640 8.110 2.390 ;
        RECT  7.850 2.110 8.080 2.390 ;
        END
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.830 0.840 9.120 2.330 ;
        END
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.400 2.040 0.720 2.360 ;
        END
    END D
    PIN CK
        DIRECTION INPUT ;
        USE clock ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.240 2.070 1.620 ;
        END
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.610 -0.280 9.200 0.280 ;
        RECT  8.330 -0.280 8.610 0.400 ;
        RECT  6.490 -0.280 8.330 0.280 ;
        RECT  6.210 -0.280 6.490 0.740 ;
        RECT  4.490 -0.280 6.210 0.280 ;
        RECT  4.330 -0.280 4.490 0.690 ;
        RECT  1.580 -0.280 4.330 0.280 ;
        RECT  1.300 -0.280 1.580 0.380 ;
        RECT  0.000 -0.280 1.300 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  8.580 3.320 9.200 3.880 ;
        RECT  7.290 3.200 8.580 3.880 ;
        RECT  6.080 3.320 7.290 3.880 ;
        RECT  5.800 3.200 6.080 3.880 ;
        RECT  3.670 3.320 5.800 3.880 ;
        RECT  3.390 2.450 3.670 3.880 ;
        RECT  2.210 3.320 3.390 3.880 ;
        RECT  1.930 3.200 2.210 3.880 ;
        RECT  0.600 3.260 1.930 3.880 ;
        RECT  0.370 3.320 0.600 3.880 ;
        RECT  0.090 3.200 0.370 3.880 ;
        RECT  0.000 3.320 0.090 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  8.640 2.600 8.920 2.880 ;
        RECT  7.010 2.680 8.640 2.880 ;
        RECT  7.670 1.670 7.730 1.950 ;
        RECT  7.670 0.450 7.710 0.670 ;
        RECT  7.650 0.450 7.670 1.950 ;
        RECT  7.510 0.450 7.650 2.520 ;
        RECT  7.430 0.450 7.510 0.670 ;
        RECT  7.490 1.410 7.510 2.520 ;
        RECT  7.370 2.240 7.490 2.520 ;
        RECT  7.010 1.030 7.350 1.310 ;
        RECT  6.850 1.030 7.010 3.160 ;
        RECT  6.290 1.900 6.850 2.060 ;
        RECT  6.260 2.940 6.850 3.160 ;
        RECT  6.470 2.500 6.690 2.780 ;
        RECT  5.730 2.500 6.470 2.660 ;
        RECT  6.010 1.780 6.290 2.060 ;
        RECT  5.570 0.790 5.730 2.880 ;
        RECT  5.450 0.790 5.570 1.070 ;
        RECT  5.190 2.720 5.570 2.880 ;
        RECT  5.130 2.310 5.410 2.560 ;
        RECT  4.970 0.790 5.190 1.830 ;
        RECT  4.910 2.720 5.190 2.990 ;
        RECT  4.750 2.310 5.130 2.470 ;
        RECT  4.370 1.670 4.970 1.830 ;
        RECT  4.590 2.310 4.750 2.940 ;
        RECT  3.990 2.780 4.590 2.940 ;
        RECT  4.370 2.340 4.430 2.620 ;
        RECT  4.150 1.670 4.370 2.620 ;
        RECT  3.850 1.170 3.990 2.940 ;
        RECT  3.830 0.760 3.850 2.940 ;
        RECT  3.690 0.760 3.830 1.330 ;
        RECT  3.090 0.760 3.690 0.920 ;
        RECT  3.510 2.010 3.670 2.290 ;
        RECT  3.410 1.080 3.530 1.300 ;
        RECT  3.410 2.010 3.510 2.170 ;
        RECT  3.250 1.080 3.410 2.170 ;
        RECT  3.230 2.010 3.250 2.170 ;
        RECT  3.070 2.010 3.230 3.020 ;
        RECT  2.910 0.760 3.090 1.660 ;
        RECT  2.770 2.860 3.070 3.020 ;
        RECT  2.750 0.760 2.910 2.460 ;
        RECT  2.490 2.860 2.770 3.080 ;
        RECT  2.550 1.910 2.750 2.460 ;
        RECT  1.100 2.300 2.550 2.460 ;
        RECT  1.220 2.860 2.490 3.020 ;
        RECT  2.230 0.860 2.390 1.960 ;
        RECT  1.760 0.860 2.230 1.080 ;
        RECT  1.740 1.800 2.230 1.960 ;
        RECT  1.460 1.800 1.740 2.130 ;
        RECT  1.040 1.800 1.460 1.960 ;
        RECT  0.940 2.620 1.220 3.020 ;
        RECT  0.880 2.180 1.100 2.460 ;
        RECT  0.880 1.720 1.040 1.960 ;
        RECT  0.240 2.620 0.940 2.780 ;
        RECT  0.620 1.720 0.880 1.880 ;
        RECT  0.400 1.340 0.620 1.880 ;
        RECT  0.240 0.900 0.370 1.180 ;
        RECT  0.080 0.900 0.240 2.790 ;
    END
END MAS91

MACRO MAS92
    CLASS CORE ;
    FOREIGN MAS92 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.310 0.440 2.320 1.560 ;
        RECT  2.120 0.440 2.310 2.330 ;
        RECT  2.080 0.440 2.120 1.560 ;
        RECT  2.080 2.080 2.120 2.330 ;
        RECT  1.120 2.120 2.080 2.280 ;
        RECT  0.960 2.120 1.120 2.470 ;
        END
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.640 1.920 1.960 ;
        RECT  1.340 1.640 1.680 1.880 ;
        END
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.520 2.600 2.120 2.780 ;
        RECT  1.280 2.440 1.520 2.780 ;
        END
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.520 0.720 1.960 ;
        END
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 1.240 1.120 1.880 ;
        END
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.920 -0.280 2.400 0.280 ;
        RECT  0.640 -0.280 0.920 0.520 ;
        RECT  0.000 -0.280 0.640 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 3.320 2.400 3.880 ;
        RECT  0.390 3.260 1.760 3.880 ;
        RECT  0.110 2.250 0.390 3.880 ;
        RECT  0.000 3.320 0.110 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  0.370 0.920 1.540 1.080 ;
        RECT  0.090 0.920 0.370 1.200 ;
    END
END MAS92

MACRO MAS93
    CLASS CORE ;
    FOREIGN MAS93 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.600 ;
    SYMMETRY x y ;
    SITE cellsite ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.770 1.030 1.990 2.760 ;
        RECT  1.680 2.440 1.770 2.760 ;
        END
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.470 1.640 2.720 2.760 ;
        RECT  2.350 1.640 2.470 1.960 ;
        RECT  2.190 0.710 2.350 1.960 ;
        RECT  1.610 0.710 2.190 0.870 ;
        RECT  1.390 0.710 1.610 1.640 ;
        END
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.480 1.520 0.910 1.960 ;
        END
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 0.440 0.320 1.740 ;
        END
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.510 -0.280 2.800 0.280 ;
        RECT  2.230 -0.280 2.510 0.340 ;
        RECT  1.370 -0.280 2.230 0.280 ;
        RECT  1.090 -0.280 1.370 0.400 ;
        RECT  0.540 -0.280 1.090 0.340 ;
        RECT  0.000 -0.280 0.540 0.280 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  2.710 3.320 2.800 3.880 ;
        RECT  2.430 3.260 2.710 3.880 ;
        RECT  1.150 3.320 2.430 3.880 ;
        RECT  0.870 3.260 1.150 3.880 ;
        RECT  0.000 3.320 0.870 3.880 ;
        END
    END VDD
    OBS
        LAYER metal1 ;
        RECT  1.520 2.940 2.190 3.160 ;
        RECT  1.230 2.940 1.520 3.100 ;
        RECT  1.070 0.980 1.230 3.100 ;
        RECT  0.790 0.980 1.070 1.140 ;
        RECT  0.310 2.940 1.070 3.100 ;
        RECT  0.510 0.860 0.790 1.140 ;
        RECT  0.150 2.030 0.310 3.100 ;
        RECT  0.090 2.030 0.150 2.830 ;
    END
END MAS93

END LIBRARY
